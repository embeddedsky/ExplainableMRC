Memristor with threshold
*.OPTIONS	POST=1	LIST ingold=2 runlvl=0
.param stime=0.5
*.param uni=unif(0.5,0.5)

* send parameters to the .control section

.csparam stime={stime}


**************MOSFET**********************************************************************
.model n12 nmos level=49 version=3.3.0 L=1.000E-05 W=1.000E-05
.model p12 pmos level=49 version=3.3.0 L=1.000E-05 W=1.000E-05

*.model n1 nmos level=49 version=3.3.0
*.model p1 pmos level=49 version=3.3.0

*.MODEL n1 NMOS level=49 version=3.3.0 W=3u L=0.35u pd=9u ad=9p ps=9u as=9p
*.MODEL p1 PMOS level=49 version=3.3.0 W=7.5u L=0.35u pd=13.5u ad=22.5p ps=13.5u as=22.5p

*.model n1 nmos level=8 version=3.2.2
*.model p1 pmos level=8 version=3.2.2

.MODEL n12 NMOS L=1.000E-05 W=1.000E-05
.MODEL p21 PMOS L=1.000E-05 W=1.000E-05

.MODEL n1 NMOS (LEVEL=49
+VERSION=3.3 CAPMOD=2 MOBMOD=1
+TOX=1E-7 NCH=1.45E17 NSUB=5.33E16 XT=8.66E-8
+VTH0=0.3 U0= 600 WINT=2.0E-7 LINT=1E-7
+NGATE=5E20 RSH=1082 JS=3.23E-8 JSW=3.23E-8 CJ=6.8E-4 MJ=0.5 PB=0.95
+CJSW=1.26E-10 MJSW=0.5 PBSW=0.95 PCLM=5
+CGSO=3.4E-10 CGDO=3.4E-10 CGBO=5.75E-10)

.MODEL p1 PMOS (LEVEL=49
+VERSION=3.3 CAPMOD=2 MOBMOD=1
+TOX=1E-7 NCH=7.12E16 NSUB=3.16E16 XT=8.66E-8
+VTH0=-0.3 U0= 376.72 WINT=2.0E-7 LINT=2.26E-7
+NGATE=5E20 RSH=1347 JS=3.51E-8 JSW=3.51E-8 CJ=5.28E-4 MJ=0.5 PB=0.94
+CJSW=1.19E-10 MJSW=0.5 PBSW=0.94
+CGSO=4.5E-10 CGDO=4.5E-10 CGBO=5.75E-10)

***************************memristor**************************************************************************************
.subckt memristor plus minus params: Ron=100 Roff=10k xini='ra' uv='1e-14/stime' p=1,

.param D=10n k={uv*Ron/pow(D,2)} a={(xini-Ron)/(Roff-xini)}

*model of memristive port
Roff plus aux {Roff}

Eres aux minus value={(Ron-Roff)/(1+a*exp(-4*k*V(q)))*I(Eres)}

*Rmem plus minus R='Roff+(Ron-Roff)/(1+a*exp(-4*k*V(q)))'
*end of the model of memristive port

*integrator model

Gx 0 Q value={i(Eres)}

Cint Q 0 1

Raux Q 0 100meg

*end of integrator model

*alternative integrator model; SDT function for PSPICE can be replaced by IDT for LTspice

*Eq Q 0 value={SDT(I(Eres))}

.ends memristor




**************reservior units-4类*********************************
***************unitrc1*********************************
.subckt unitrc1 in out params: ra=0.14 tb=0.03
xmen 2 121 memristor xini='ra'
vtemp2 121 1 dc 0
Mp1 2 cpminus in in p1
Mn1 1 cppulse out out n1
Mn2 2 cpminus out out n1
Mp2 1 cppulse in in p1
vcp41 cppulse 0 DC 0 PULSE(0 5 0 0 0 'tb*stime' 'tb*2*stime')
vcp42 cpminus 0 DC 0 PULSE(5 0 0 0 0 'tb*stime' 'tb*2*stime')
*vtemp1 out1 out dc 0
*xs1 out2 0 out myswitch
.ends


***************unitrc3（大阻值相当于断路）*********************************
.subckt unitrc2 in out
R1 in out 1e+12
.ends

***********input voltage*****************
*vcp 100 0 sin(2.5 2.5 '10/stime' 0 0 0)
*vcp 100 0 sin(4.5 4.5 '20/stime' '0.5*stime' 0 0)
.subckt filesource1 1 2
a1 %vd([1 2]) filesrc1
.model filesrc1 filesource (file="signal1.m" amploffset=[0] amplscale=[1]
+ timeoffset=0 timescale=1
+ timerelative=false amplstep=false)
.ends

.subckt filesource2 1 2
a1 %vd([1 2]) filesrc2
.model filesrc2 filesource (file="signal2.m" amploffset=[0] amplscale=[1]
+ timeoffset=0 timescale=1
+ timerelative=false amplstep=false)
.ends

.subckt filesource3 1 2
a1 %vd([1 2]) filesrc3
.model filesrc3 filesource (file="signal3.m" amploffset=[0] amplscale=[1]
+ timeoffset=0 timescale=1
+ timerelative=false amplstep=false)
.ends

.subckt filesource4 1 2
a1 %vd([1 2]) filesrc4
.model filesrc4 filesource (file="signal1.m" amploffset=[0] amplscale=[1]
+ timeoffset=0 timescale=1
+ timerelative=false amplstep=false)
.ends

.subckt filesource5 1 2
a1 %vd([1 2]) filesrc5
.model filesrc5 filesource (file="signal2.m" amploffset=[0] amplscale=[1]
+ timeoffset=0 timescale=1
+ timerelative=false amplstep=false)
.ends

.subckt filesource6 1 2
a1 %vd([1 2]) filesrc6
.model filesrc6 filesource (file="signal3.m" amploffset=[0] amplscale=[1]
+ timeoffset=0 timescale=1
+ timerelative=false amplstep=false)
.ends

.subckt filesource7 1 2
a1 %vd([1 2]) filesrc7
.model filesrc7 filesource (file="signal1.m" amploffset=[0] amplscale=[1]
+ timeoffset=0 timescale=1
+ timerelative=false amplstep=false)
.ends

.subckt filesource8 1 2
a1 %vd([1 2]) filesrc8
.model filesrc8 filesource (file="signal2.m" amploffset=[0] amplscale=[1]
+ timeoffset=0 timescale=1
+ timerelative=false amplstep=false)
.ends

.subckt filesource9 1 2
a1 %vd([1 2]) filesrc9
.model filesrc9 filesource (file="signal3.m" amploffset=[0] amplscale=[1]
+ timeoffset=0 timescale=1
+ timerelative=false amplstep=false)
.ends

X1 100 0 filesource1
X2 101 0 filesource2
X3 102 0 filesource3
X4 103 0 filesource4
X5 104 0 filesource5
X6 105 0 filesource6
X7 106 0 filesource7
X8 107 0 filesource8
X9 108 0 filesource9
***********target voltage*****************
*vtarget1 vt1 0 DC 0 PULSE(0 0.001 0 0 0 'stime/20' 'stime/10')
*vtarget2 vt2 0 DC 0 PULSE(0 0.001 0  'stime/20' 0 'stime/999' 'stime/10')
*vtarget3 vt3 0 DC 0 sin(0.0005 0.0005 '20/stime' 0 0 0)

.subckt filesource10 1 2
a1 %vd([1 2]) filesrc10
.model filesrc10 filesource (file="output.m" amploffset=[0] amplscale=[1]
+ timeoffset=0 timescale=1
+ timerelative=false amplstep=false)
.ends

xtarget1 vt1 0 filesource10
**************input layer***********
*xunitin1 1 2 unitin ta=0.199
*xopein 2 5 ope
*Rin1 1 5 1k
***********reservior input voltage (演化下面out_gain这个参数-1到1之间)*****************
*vp1 112 0 DC 0 PULSE(1 0 0 0 0 'stime' 'stime')
*a2 [5 112] 113 sigmulta2
*.model sigmulta2 mult(in_offset=[0 0]
*+ in_gain=[1.0 1.0] out_gain=1 out_offset=0)

************待生成reservior*(必须包含节点113)(6-26)*********************************
*************随机选择reservior中的一个节点接输入和地***********


vtemprc1 100 21 dc 0
vtemprc2 101 13 dc 0
vtemprc3 102 1 dc 0
vtemprc4 103 48 dc 0
vtemprc5 104 4 dc 0
vtemprc6 105 8 dc 0
vtemprc7 106 28 dc 0
vtemprc8 107 11 dc 0
vtemprc9 108 23 dc 0
vtemprc10  39 0 dc 0
xunit1-1  1  1  unitrc1  ra=6383.76  tb=0.26
xunit1-2  1  2  unitrc1  ra=6325.17  tb=0.41
xunit1-4  1  4  unitrc1  ra=7986.39  tb=0.19
xunit1-6  1  6  unitrc1  ra=2058.48  tb=0.35
xunit1-8  1  8  unitrc1  ra=2173.10  tb=0.05
xunit1-9  1  9  unitrc1  ra=3663.51  tb=0.21
xunit1-10  1  10  unitrc1  ra=6279.56  tb=0.15
xunit1-14  1  14  unitrc1  ra=1853.74  tb=0.39
xunit1-15  1  15  unitrc1  ra=9982.65  tb=0.23
xunit1-16  1  16  unitrc1  ra=3317.93  tb=0.13
xunit1-17  1  17  unitrc1  ra=8276.86  tb=0.30
xunit1-18  1  18  unitrc1  ra=8330.58  tb=0.22
xunit1-21  1  21  unitrc1  ra=7548.66  tb=0.40
xunit1-22  1  22  unitrc1  ra=6905.26  tb=0.17
xunit1-23  1  23  unitrc1  ra=4931.23  tb=0.22
xunit1-24  1  24  unitrc1  ra=1694.38  tb=0.41
xunit1-25  1  25  unitrc1  ra=8294.53  tb=0.25
xunit1-26  1  26  unitrc1  ra=8747.66  tb=0.49
xunit1-27  1  27  unitrc1  ra=1500.27  tb=0.08
xunit1-29  1  29  unitrc1  ra=2043.43  tb=0.45
xunit1-32  1  32  unitrc1  ra=4698.16  tb=0.03
xunit1-34  1  34  unitrc1  ra=2525.33  tb=0.35
xunit1-35  1  35  unitrc1  ra=305.57  tb=0.07
xunit1-42  1  42  unitrc1  ra=4061.78  tb=0.19
xunit1-45  1  45  unitrc1  ra=4519.64  tb=0.24
xunit1-46  1  46  unitrc1  ra=2179.21  tb=0.04

xunit2-1  2  1  unitrc1  ra=8454.72  tb=0.09
xunit2-3  2  3  unitrc1  ra=3248.39  tb=0.20
xunit2-8  2  8  unitrc1  ra=2297.76  tb=0.50
xunit2-12  2  12  unitrc1  ra=2005.72  tb=0.18
xunit2-13  2  13  unitrc1  ra=316.63  tb=0.12
xunit2-14  2  14  unitrc1  ra=5377.89  tb=0.10
xunit2-15  2  15  unitrc1  ra=9613.83  tb=0.15
xunit2-16  2  16  unitrc1  ra=6959.19  tb=0.18
xunit2-17  2  17  unitrc1  ra=8410.07  tb=0.50
xunit2-18  2  18  unitrc1  ra=9120.85  tb=0.37
xunit2-19  2  19  unitrc1  ra=7786.26  tb=0.30
xunit2-20  2  20  unitrc1  ra=3738.96  tb=0.34
xunit2-22  2  22  unitrc1  ra=6208.83  tb=0.35
xunit2-23  2  23  unitrc1  ra=4445.05  tb=0.28
xunit2-24  2  24  unitrc1  ra=1637.95  tb=0.29
xunit2-27  2  27  unitrc1  ra=3320.00  tb=0.48
xunit2-32  2  32  unitrc1  ra=3856.00  tb=0.00
xunit2-36  2  36  unitrc1  ra=4990.51  tb=0.24
xunit2-39  2  39  unitrc1  ra=9943.29  tb=0.38
xunit2-40  2  40  unitrc1  ra=2598.66  tb=0.32
xunit2-41  2  41  unitrc1  ra=4358.08  tb=0.43
xunit2-43  2  43  unitrc1  ra=6600.96  tb=0.01
xunit2-44  2  44  unitrc1  ra=7904.19  tb=0.13
xunit2-45  2  45  unitrc1  ra=6317.24  tb=0.36
xunit2-46  2  46  unitrc1  ra=4116.29  tb=0.41
xunit2-47  2  47  unitrc1  ra=6210.64  tb=0.18
xunit2-48  2  48  unitrc1  ra=673.18  tb=0.10

xunit3-2  3  2  unitrc1  ra=5770.45  tb=0.37
xunit3-3  3  3  unitrc1  ra=7072.86  tb=0.37
xunit3-4  3  4  unitrc1  ra=2679.23  tb=0.00
xunit3-6  3  6  unitrc1  ra=3590.44  tb=0.32
xunit3-7  3  7  unitrc1  ra=9412.52  tb=0.08
xunit3-8  3  8  unitrc1  ra=5378.42  tb=0.23
xunit3-11  3  11  unitrc1  ra=832.19  tb=0.15
xunit3-12  3  12  unitrc1  ra=4333.41  tb=0.49
xunit3-15  3  15  unitrc1  ra=410.54  tb=0.39
xunit3-16  3  16  unitrc1  ra=3456.86  tb=0.18
xunit3-18  3  18  unitrc1  ra=3836.13  tb=0.22
xunit3-20  3  20  unitrc1  ra=6699.62  tb=0.31
xunit3-22  3  22  unitrc1  ra=1733.38  tb=0.32
xunit3-23  3  23  unitrc1  ra=5680.87  tb=0.22
xunit3-25  3  25  unitrc1  ra=8207.55  tb=0.33
xunit3-26  3  26  unitrc1  ra=5074.03  tb=0.49
xunit3-27  3  27  unitrc1  ra=9584.14  tb=0.14
xunit3-32  3  32  unitrc1  ra=5276.00  tb=0.40
xunit3-36  3  36  unitrc1  ra=3858.92  tb=0.14
xunit3-37  3  37  unitrc1  ra=5892.31  tb=0.47
xunit3-39  3  39  unitrc1  ra=7981.20  tb=0.06
xunit3-43  3  43  unitrc1  ra=5673.27  tb=0.29
xunit3-45  3  45  unitrc1  ra=1864.28  tb=0.44
xunit3-48  3  48  unitrc1  ra=3953.70  tb=0.13
xunit3-49  3  49  unitrc1  ra=5085.58  tb=0.24
xunit3-50  3  50  unitrc1  ra=782.84  tb=0.06

xunit4-1  4  1  unitrc1  ra=2020.83  tb=0.27
xunit4-3  4  3  unitrc1  ra=1976.48  tb=0.01
xunit4-4  4  4  unitrc1  ra=2882.75  tb=0.17
xunit4-5  4  5  unitrc1  ra=9345.15  tb=0.12
xunit4-7  4  7  unitrc1  ra=2535.95  tb=0.39
xunit4-8  4  8  unitrc1  ra=4046.51  tb=0.45
xunit4-9  4  9  unitrc1  ra=448.97  tb=0.38
xunit4-14  4  14  unitrc1  ra=6124.20  tb=0.09
xunit4-15  4  15  unitrc1  ra=1178.61  tb=0.17
xunit4-16  4  16  unitrc1  ra=500.15  tb=0.19
xunit4-18  4  18  unitrc1  ra=6545.71  tb=0.21
xunit4-19  4  19  unitrc1  ra=6365.49  tb=0.32
xunit4-20  4  20  unitrc1  ra=807.78  tb=0.34
xunit4-21  4  21  unitrc1  ra=3505.45  tb=0.16
xunit4-24  4  24  unitrc1  ra=5493.13  tb=0.14
xunit4-25  4  25  unitrc1  ra=1964.26  tb=0.11
xunit4-26  4  26  unitrc1  ra=2781.86  tb=0.43
xunit4-27  4  27  unitrc1  ra=3840.66  tb=0.08
xunit4-28  4  28  unitrc1  ra=8989.84  tb=0.03
xunit4-29  4  29  unitrc1  ra=7456.39  tb=0.24
xunit4-33  4  33  unitrc1  ra=3569.37  tb=0.29
xunit4-34  4  34  unitrc1  ra=1335.94  tb=0.16
xunit4-35  4  35  unitrc1  ra=4072.00  tb=0.48
xunit4-36  4  36  unitrc1  ra=8787.59  tb=0.14
xunit4-37  4  37  unitrc1  ra=8709.14  tb=0.04
xunit4-38  4  38  unitrc1  ra=4219.53  tb=0.36
xunit4-39  4  39  unitrc1  ra=2793.97  tb=0.11
xunit4-41  4  41  unitrc1  ra=4422.97  tb=0.14
xunit4-42  4  42  unitrc1  ra=4279.63  tb=0.15
xunit4-47  4  47  unitrc1  ra=4034.72  tb=0.06
xunit4-49  4  49  unitrc1  ra=6556.42  tb=0.36
xunit4-50  4  50  unitrc1  ra=2454.08  tb=0.28

xunit5-1  5  1  unitrc1  ra=844.83  tb=0.04
xunit5-3  5  3  unitrc1  ra=4635.80  tb=0.12
xunit5-5  5  5  unitrc1  ra=9609.57  tb=0.40
xunit5-6  5  6  unitrc1  ra=9618.94  tb=0.15
xunit5-8  5  8  unitrc1  ra=2779.11  tb=0.43
xunit5-9  5  9  unitrc1  ra=3945.77  tb=0.11
xunit5-12  5  12  unitrc1  ra=9034.16  tb=0.19
xunit5-13  5  13  unitrc1  ra=5267.29  tb=0.18
xunit5-14  5  14  unitrc1  ra=2193.40  tb=0.43
xunit5-16  5  16  unitrc1  ra=7900.84  tb=0.10
xunit5-17  5  17  unitrc1  ra=9864.62  tb=0.22
xunit5-18  5  18  unitrc1  ra=6086.12  tb=0.11
xunit5-19  5  19  unitrc1  ra=5806.04  tb=0.15
xunit5-20  5  20  unitrc1  ra=7848.21  tb=0.08
xunit5-21  5  21  unitrc1  ra=4472.35  tb=0.14
xunit5-23  5  23  unitrc1  ra=4599.71  tb=0.11
xunit5-27  5  27  unitrc1  ra=5424.35  tb=0.37
xunit5-28  5  28  unitrc1  ra=6074.26  tb=0.46
xunit5-29  5  29  unitrc1  ra=348.66  tb=0.34
xunit5-31  5  31  unitrc1  ra=5413.29  tb=0.24
xunit5-32  5  32  unitrc1  ra=2206.72  tb=0.20
xunit5-33  5  33  unitrc1  ra=1018.06  tb=0.46
xunit5-37  5  37  unitrc1  ra=5777.31  tb=0.27
xunit5-39  5  39  unitrc1  ra=3959.67  tb=0.22
xunit5-43  5  43  unitrc1  ra=6399.41  tb=0.30
xunit5-44  5  44  unitrc1  ra=4830.54  tb=0.08
xunit5-45  5  45  unitrc1  ra=1956.41  tb=0.14
xunit5-47  5  47  unitrc1  ra=1838.89  tb=0.17
xunit5-49  5  49  unitrc1  ra=5852.01  tb=0.46
xunit5-50  5  50  unitrc1  ra=3836.31  tb=0.21

xunit6-1  6  1  unitrc1  ra=4361.17  tb=0.31
xunit6-2  6  2  unitrc1  ra=1225.17  tb=0.28
xunit6-3  6  3  unitrc1  ra=3477.85  tb=0.02
xunit6-4  6  4  unitrc1  ra=2042.93  tb=0.49
xunit6-5  6  5  unitrc1  ra=2775.92  tb=0.38
xunit6-7  6  7  unitrc1  ra=3185.70  tb=0.41
xunit6-8  6  8  unitrc1  ra=2602.30  tb=0.31
xunit6-10  6  10  unitrc1  ra=4142.22  tb=0.23
xunit6-11  6  11  unitrc1  ra=7896.59  tb=0.06
xunit6-12  6  12  unitrc1  ra=3262.57  tb=0.40
xunit6-13  6  13  unitrc1  ra=7777.33  tb=0.11
xunit6-14  6  14  unitrc1  ra=613.28  tb=0.02
xunit6-15  6  15  unitrc1  ra=2471.67  tb=0.25
xunit6-16  6  16  unitrc1  ra=1757.82  tb=0.32
xunit6-17  6  17  unitrc1  ra=7259.77  tb=0.29
xunit6-18  6  18  unitrc1  ra=8219.14  tb=0.05
xunit6-21  6  21  unitrc1  ra=416.97  tb=0.16
xunit6-22  6  22  unitrc1  ra=1886.39  tb=0.16
xunit6-26  6  26  unitrc1  ra=9177.22  tb=0.24
xunit6-28  6  28  unitrc1  ra=1464.43  tb=0.14
xunit6-29  6  29  unitrc1  ra=4980.52  tb=0.36
xunit6-31  6  31  unitrc1  ra=3502.89  tb=0.22
xunit6-33  6  33  unitrc1  ra=501.80  tb=0.04
xunit6-34  6  34  unitrc1  ra=5757.22  tb=0.30
xunit6-37  6  37  unitrc1  ra=4850.07  tb=0.40
xunit6-38  6  38  unitrc1  ra=3360.98  tb=0.14
xunit6-39  6  39  unitrc1  ra=193.57  tb=0.37
xunit6-42  6  42  unitrc1  ra=8964.89  tb=0.21
xunit6-45  6  45  unitrc1  ra=1657.83  tb=0.38
xunit6-46  6  46  unitrc1  ra=4707.85  tb=0.16
xunit6-47  6  47  unitrc1  ra=9733.85  tb=0.35
xunit6-48  6  48  unitrc1  ra=2852.43  tb=0.23
xunit6-49  6  49  unitrc1  ra=6308.80  tb=0.44

xunit7-4  7  4  unitrc1  ra=4732.17  tb=0.04
xunit7-5  7  5  unitrc1  ra=556.25  tb=0.03
xunit7-6  7  6  unitrc1  ra=2458.92  tb=0.32
xunit7-8  7  8  unitrc1  ra=8348.91  tb=0.37
xunit7-9  7  9  unitrc1  ra=1717.15  tb=0.39
xunit7-10  7  10  unitrc1  ra=3614.99  tb=0.09
xunit7-13  7  13  unitrc1  ra=2705.59  tb=0.37
xunit7-14  7  14  unitrc1  ra=7122.73  tb=0.37
xunit7-15  7  15  unitrc1  ra=8162.74  tb=0.32
xunit7-16  7  16  unitrc1  ra=455.44  tb=0.48
xunit7-17  7  17  unitrc1  ra=8527.68  tb=0.45
xunit7-19  7  19  unitrc1  ra=4988.46  tb=0.34
xunit7-21  7  21  unitrc1  ra=4836.12  tb=0.42
xunit7-24  7  24  unitrc1  ra=3661.52  tb=0.39
xunit7-25  7  25  unitrc1  ra=8898.18  tb=0.30
xunit7-26  7  26  unitrc1  ra=2479.38  tb=0.34
xunit7-27  7  27  unitrc1  ra=2685.50  tb=0.10
xunit7-32  7  32  unitrc1  ra=8810.44  tb=0.29
xunit7-33  7  33  unitrc1  ra=2704.85  tb=0.32
xunit7-34  7  34  unitrc1  ra=3108.80  tb=0.27
xunit7-35  7  35  unitrc1  ra=6939.10  tb=0.22
xunit7-36  7  36  unitrc1  ra=152.60  tb=0.37
xunit7-40  7  40  unitrc1  ra=5282.79  tb=0.48
xunit7-42  7  42  unitrc1  ra=8482.62  tb=0.44
xunit7-44  7  44  unitrc1  ra=5063.30  tb=0.09
xunit7-45  7  45  unitrc1  ra=4125.29  tb=0.42
xunit7-46  7  46  unitrc1  ra=6401.14  tb=0.24
xunit7-47  7  47  unitrc1  ra=8149.57  tb=0.03
xunit7-48  7  48  unitrc1  ra=4062.62  tb=0.17
xunit7-50  7  50  unitrc1  ra=4826.78  tb=0.05

xunit8-3  8  3  unitrc1  ra=6761.18  tb=0.49
xunit8-5  8  5  unitrc1  ra=8788.63  tb=0.04
xunit8-6  8  6  unitrc1  ra=3041.27  tb=0.27
xunit8-8  8  8  unitrc1  ra=352.73  tb=0.47
xunit8-9  8  9  unitrc1  ra=150.16  tb=0.10
xunit8-10  8  10  unitrc1  ra=1730.90  tb=0.30
xunit8-11  8  11  unitrc1  ra=7943.92  tb=0.38
xunit8-13  8  13  unitrc1  ra=742.88  tb=0.46
xunit8-15  8  15  unitrc1  ra=1749.41  tb=0.17
xunit8-16  8  16  unitrc1  ra=8856.15  tb=0.29
xunit8-17  8  17  unitrc1  ra=699.86  tb=0.14
xunit8-18  8  18  unitrc1  ra=7579.63  tb=0.29
xunit8-20  8  20  unitrc1  ra=4398.01  tb=0.40
xunit8-22  8  22  unitrc1  ra=6217.31  tb=0.42
xunit8-24  8  24  unitrc1  ra=6948.47  tb=0.19
xunit8-25  8  25  unitrc1  ra=2133.60  tb=0.10
xunit8-29  8  29  unitrc1  ra=2580.30  tb=0.17
xunit8-30  8  30  unitrc1  ra=2942.71  tb=0.39
xunit8-31  8  31  unitrc1  ra=762.02  tb=0.23
xunit8-32  8  32  unitrc1  ra=6235.92  tb=0.46
xunit8-37  8  37  unitrc1  ra=5515.28  tb=0.08
xunit8-40  8  40  unitrc1  ra=4227.40  tb=0.03
xunit8-42  8  42  unitrc1  ra=195.00  tb=0.40
xunit8-43  8  43  unitrc1  ra=2363.07  tb=0.20
xunit8-45  8  45  unitrc1  ra=4694.27  tb=0.10
xunit8-48  8  48  unitrc1  ra=4467.83  tb=0.24
xunit8-49  8  49  unitrc1  ra=9642.88  tb=0.07

xunit9-1  9  1  unitrc1  ra=6775.66  tb=0.48
xunit9-2  9  2  unitrc1  ra=9208.10  tb=0.37
xunit9-4  9  4  unitrc1  ra=8092.85  tb=0.49
xunit9-5  9  5  unitrc1  ra=9093.97  tb=0.19
xunit9-6  9  6  unitrc1  ra=2561.61  tb=0.34
xunit9-8  9  8  unitrc1  ra=3847.96  tb=0.36
xunit9-9  9  9  unitrc1  ra=8169.50  tb=0.14
xunit9-10  9  10  unitrc1  ra=8019.50  tb=0.13
xunit9-11  9  11  unitrc1  ra=3704.93  tb=0.36
xunit9-12  9  12  unitrc1  ra=6109.11  tb=0.16
xunit9-13  9  13  unitrc1  ra=3777.40  tb=0.13
xunit9-16  9  16  unitrc1  ra=2387.29  tb=0.44
xunit9-17  9  17  unitrc1  ra=8675.62  tb=0.08
xunit9-18  9  18  unitrc1  ra=517.68  tb=0.13
xunit9-19  9  19  unitrc1  ra=3993.91  tb=0.31
xunit9-21  9  21  unitrc1  ra=3732.66  tb=0.07
xunit9-22  9  22  unitrc1  ra=5574.63  tb=0.47
xunit9-23  9  23  unitrc1  ra=7535.76  tb=0.08
xunit9-24  9  24  unitrc1  ra=8560.33  tb=0.37
xunit9-25  9  25  unitrc1  ra=5231.55  tb=0.45
xunit9-27  9  27  unitrc1  ra=1699.86  tb=0.13
xunit9-34  9  34  unitrc1  ra=6844.57  tb=0.15
xunit9-35  9  35  unitrc1  ra=6223.32  tb=0.49
xunit9-36  9  36  unitrc1  ra=7844.01  tb=0.20
xunit9-37  9  37  unitrc1  ra=3261.64  tb=0.38
xunit9-38  9  38  unitrc1  ra=4428.81  tb=0.47
xunit9-39  9  39  unitrc1  ra=4046.11  tb=0.35
xunit9-40  9  40  unitrc1  ra=4381.20  tb=0.15
xunit9-41  9  41  unitrc1  ra=591.82  tb=0.20
xunit9-45  9  45  unitrc1  ra=1715.72  tb=0.08
xunit9-46  9  46  unitrc1  ra=3845.81  tb=0.38
xunit9-47  9  47  unitrc1  ra=3452.34  tb=0.03
xunit9-49  9  49  unitrc1  ra=6559.87  tb=0.47

xunit10-1  10  1  unitrc1  ra=272.67  tb=0.28
xunit10-4  10  4  unitrc1  ra=8253.12  tb=0.44
xunit10-7  10  7  unitrc1  ra=6850.57  tb=0.14
xunit10-8  10  8  unitrc1  ra=4225.32  tb=0.29
xunit10-9  10  9  unitrc1  ra=5013.43  tb=0.32
xunit10-10  10  10  unitrc1  ra=6114.43  tb=0.19
xunit10-11  10  11  unitrc1  ra=9775.08  tb=0.08
xunit10-12  10  12  unitrc1  ra=1992.99  tb=0.27
xunit10-14  10  14  unitrc1  ra=5284.04  tb=0.19
xunit10-15  10  15  unitrc1  ra=2052.74  tb=0.25
xunit10-16  10  16  unitrc1  ra=7119.17  tb=0.38
xunit10-18  10  18  unitrc1  ra=8182.41  tb=0.34
xunit10-19  10  19  unitrc1  ra=9254.65  tb=0.23
xunit10-21  10  21  unitrc1  ra=3800.34  tb=0.02
xunit10-23  10  23  unitrc1  ra=4238.63  tb=0.28
xunit10-26  10  26  unitrc1  ra=5430.87  tb=0.05
xunit10-28  10  28  unitrc1  ra=161.56  tb=0.27
xunit10-29  10  29  unitrc1  ra=3709.14  tb=0.13
xunit10-30  10  30  unitrc1  ra=8758.01  tb=0.12
xunit10-32  10  32  unitrc1  ra=4674.47  tb=0.19
xunit10-33  10  33  unitrc1  ra=8021.42  tb=0.25
xunit10-34  10  34  unitrc1  ra=371.23  tb=0.20
xunit10-35  10  35  unitrc1  ra=8051.67  tb=0.07
xunit10-36  10  36  unitrc1  ra=4042.86  tb=0.19
xunit10-37  10  37  unitrc1  ra=2678.47  tb=0.45
xunit10-38  10  38  unitrc1  ra=414.27  tb=0.26
xunit10-39  10  39  unitrc1  ra=3970.41  tb=0.26
xunit10-41  10  41  unitrc1  ra=3383.06  tb=0.06
xunit10-42  10  42  unitrc1  ra=4052.73  tb=0.41
xunit10-43  10  43  unitrc1  ra=1438.85  tb=0.15
xunit10-45  10  45  unitrc1  ra=7799.25  tb=0.36
xunit10-46  10  46  unitrc1  ra=2744.63  tb=0.41
xunit10-47  10  47  unitrc1  ra=3471.04  tb=0.14
xunit10-49  10  49  unitrc1  ra=7024.23  tb=0.38
xunit10-50  10  50  unitrc1  ra=8818.13  tb=0.33

xunit11-1  11  1  unitrc1  ra=3293.28  tb=0.30
xunit11-3  11  3  unitrc1  ra=2187.12  tb=0.46
xunit11-5  11  5  unitrc1  ra=832.83  tb=0.43
xunit11-6  11  6  unitrc1  ra=6816.90  tb=0.05
xunit11-7  11  7  unitrc1  ra=1922.19  tb=0.22
xunit11-8  11  8  unitrc1  ra=1388.29  tb=0.06
xunit11-9  11  9  unitrc1  ra=1254.88  tb=0.26
xunit11-10  11  10  unitrc1  ra=2949.15  tb=0.25
xunit11-12  11  12  unitrc1  ra=5835.92  tb=0.08
xunit11-13  11  13  unitrc1  ra=2517.63  tb=0.12
xunit11-15  11  15  unitrc1  ra=2834.63  tb=0.32
xunit11-16  11  16  unitrc1  ra=8002.21  tb=0.42
xunit11-18  11  18  unitrc1  ra=5413.96  tb=0.47
xunit11-19  11  19  unitrc1  ra=7667.56  tb=0.36
xunit11-20  11  20  unitrc1  ra=3829.79  tb=0.12
xunit11-21  11  21  unitrc1  ra=908.00  tb=0.24
xunit11-22  11  22  unitrc1  ra=585.33  tb=0.49
xunit11-23  11  23  unitrc1  ra=3015.04  tb=0.50
xunit11-24  11  24  unitrc1  ra=5075.75  tb=0.07
xunit11-25  11  25  unitrc1  ra=1693.40  tb=0.12
xunit11-27  11  27  unitrc1  ra=494.38  tb=0.05
xunit11-32  11  32  unitrc1  ra=4900.37  tb=0.40
xunit11-34  11  34  unitrc1  ra=5093.39  tb=0.24
xunit11-35  11  35  unitrc1  ra=6996.56  tb=0.43
xunit11-36  11  36  unitrc1  ra=676.48  tb=0.17
xunit11-37  11  37  unitrc1  ra=5056.59  tb=0.34
xunit11-38  11  38  unitrc1  ra=5288.82  tb=0.05
xunit11-39  11  39  unitrc1  ra=5937.73  tb=0.47
xunit11-40  11  40  unitrc1  ra=5804.79  tb=0.36
xunit11-43  11  43  unitrc1  ra=5057.50  tb=0.16
xunit11-45  11  45  unitrc1  ra=6169.39  tb=0.19
xunit11-47  11  47  unitrc1  ra=4380.31  tb=0.43
xunit11-48  11  48  unitrc1  ra=5714.28  tb=0.00
xunit11-49  11  49  unitrc1  ra=3407.36  tb=0.43

xunit12-1  12  1  unitrc1  ra=5870.86  tb=0.49
xunit12-2  12  2  unitrc1  ra=4987.98  tb=0.24
xunit12-4  12  4  unitrc1  ra=7198.54  tb=0.03
xunit12-5  12  5  unitrc1  ra=2498.70  tb=0.17
xunit12-7  12  7  unitrc1  ra=1978.65  tb=0.35
xunit12-9  12  9  unitrc1  ra=317.61  tb=0.26
xunit12-11  12  11  unitrc1  ra=5050.67  tb=0.07
xunit12-13  12  13  unitrc1  ra=8210.63  tb=0.17
xunit12-14  12  14  unitrc1  ra=3108.99  tb=0.13
xunit12-15  12  15  unitrc1  ra=3223.96  tb=0.19
xunit12-16  12  16  unitrc1  ra=2937.10  tb=0.37
xunit12-17  12  17  unitrc1  ra=5410.95  tb=0.28
xunit12-18  12  18  unitrc1  ra=4177.14  tb=0.03
xunit12-20  12  20  unitrc1  ra=1824.95  tb=0.23
xunit12-24  12  24  unitrc1  ra=2984.99  tb=0.42
xunit12-26  12  26  unitrc1  ra=2150.75  tb=0.36
xunit12-28  12  28  unitrc1  ra=5674.76  tb=0.31
xunit12-29  12  29  unitrc1  ra=3578.33  tb=0.24
xunit12-32  12  32  unitrc1  ra=4814.01  tb=0.21
xunit12-33  12  33  unitrc1  ra=7691.86  tb=0.47
xunit12-34  12  34  unitrc1  ra=5945.02  tb=0.25
xunit12-35  12  35  unitrc1  ra=6095.82  tb=0.20
xunit12-37  12  37  unitrc1  ra=1934.79  tb=0.26
xunit12-38  12  38  unitrc1  ra=5384.94  tb=0.38
xunit12-42  12  42  unitrc1  ra=2720.03  tb=0.43
xunit12-44  12  44  unitrc1  ra=3333.32  tb=0.03
xunit12-45  12  45  unitrc1  ra=3443.65  tb=0.34
xunit12-46  12  46  unitrc1  ra=4459.56  tb=0.05
xunit12-47  12  47  unitrc1  ra=7799.03  tb=0.34
xunit12-49  12  49  unitrc1  ra=1682.37  tb=0.22

xunit13-1  13  1  unitrc1  ra=2216.29  tb=0.47
xunit13-6  13  6  unitrc1  ra=6918.68  tb=0.33
xunit13-7  13  7  unitrc1  ra=659.23  tb=0.37
xunit13-10  13  10  unitrc1  ra=2999.72  tb=0.30
xunit13-11  13  11  unitrc1  ra=3855.62  tb=0.17
xunit13-12  13  12  unitrc1  ra=6550.72  tb=0.08
xunit13-13  13  13  unitrc1  ra=3967.19  tb=0.29
xunit13-14  13  14  unitrc1  ra=7254.96  tb=0.17
xunit13-15  13  15  unitrc1  ra=9986.07  tb=0.20
xunit13-18  13  18  unitrc1  ra=4059.40  tb=0.34
xunit13-20  13  20  unitrc1  ra=3298.37  tb=0.19
xunit13-21  13  21  unitrc1  ra=7337.74  tb=0.36
xunit13-22  13  22  unitrc1  ra=7156.46  tb=0.12
xunit13-23  13  23  unitrc1  ra=3683.49  tb=0.34
xunit13-24  13  24  unitrc1  ra=1791.92  tb=0.39
xunit13-30  13  30  unitrc1  ra=9849.05  tb=0.02
xunit13-31  13  31  unitrc1  ra=7137.47  tb=0.04
xunit13-33  13  33  unitrc1  ra=8992.00  tb=0.23
xunit13-36  13  36  unitrc1  ra=5049.06  tb=0.08
xunit13-37  13  37  unitrc1  ra=2885.77  tb=0.11
xunit13-42  13  42  unitrc1  ra=7734.89  tb=0.05
xunit13-43  13  43  unitrc1  ra=6284.96  tb=0.36
xunit13-44  13  44  unitrc1  ra=4195.98  tb=0.14
xunit13-47  13  47  unitrc1  ra=4007.79  tb=0.00
xunit13-48  13  48  unitrc1  ra=8374.20  tb=0.42
xunit13-50  13  50  unitrc1  ra=7781.64  tb=0.26

xunit14-1  14  1  unitrc1  ra=1417.08  tb=0.15
xunit14-2  14  2  unitrc1  ra=7643.50  tb=0.26
xunit14-3  14  3  unitrc1  ra=1710.49  tb=0.10
xunit14-4  14  4  unitrc1  ra=2255.72  tb=0.30
xunit14-7  14  7  unitrc1  ra=7668.65  tb=0.38
xunit14-8  14  8  unitrc1  ra=2957.15  tb=0.12
xunit14-12  14  12  unitrc1  ra=5547.26  tb=0.42
xunit14-13  14  13  unitrc1  ra=1907.97  tb=0.42
xunit14-14  14  14  unitrc1  ra=4588.46  tb=0.10
xunit14-15  14  15  unitrc1  ra=3724.69  tb=0.32
xunit14-16  14  16  unitrc1  ra=1446.98  tb=0.25
xunit14-20  14  20  unitrc1  ra=3677.29  tb=0.21
xunit14-21  14  21  unitrc1  ra=958.17  tb=0.16
xunit14-22  14  22  unitrc1  ra=1259.33  tb=0.45
xunit14-23  14  23  unitrc1  ra=4595.57  tb=0.36
xunit14-25  14  25  unitrc1  ra=4590.89  tb=0.32
xunit14-26  14  26  unitrc1  ra=6818.24  tb=0.28
xunit14-30  14  30  unitrc1  ra=3248.64  tb=0.00
xunit14-31  14  31  unitrc1  ra=3420.47  tb=0.36
xunit14-32  14  32  unitrc1  ra=8673.91  tb=0.29
xunit14-35  14  35  unitrc1  ra=8158.54  tb=0.45
xunit14-36  14  36  unitrc1  ra=9063.34  tb=0.06
xunit14-38  14  38  unitrc1  ra=2877.79  tb=0.28
xunit14-39  14  39  unitrc1  ra=6219.96  tb=0.14
xunit14-40  14  40  unitrc1  ra=1997.60  tb=0.18
xunit14-42  14  42  unitrc1  ra=4807.93  tb=0.17
xunit14-43  14  43  unitrc1  ra=2220.79  tb=0.33
xunit14-44  14  44  unitrc1  ra=2573.35  tb=0.38
xunit14-45  14  45  unitrc1  ra=888.65  tb=0.48
xunit14-46  14  46  unitrc1  ra=6566.97  tb=0.09
xunit14-48  14  48  unitrc1  ra=5654.02  tb=0.02
xunit14-49  14  49  unitrc1  ra=5702.06  tb=0.29

xunit15-1  15  1  unitrc1  ra=8045.97  tb=0.35
xunit15-2  15  2  unitrc1  ra=4279.82  tb=0.46
xunit15-3  15  3  unitrc1  ra=5321.92  tb=0.19
xunit15-5  15  5  unitrc1  ra=1826.58  tb=0.25
xunit15-9  15  9  unitrc1  ra=4495.65  tb=0.19
xunit15-11  15  11  unitrc1  ra=1845.55  tb=0.33
xunit15-13  15  13  unitrc1  ra=5841.15  tb=0.37
xunit15-14  15  14  unitrc1  ra=8126.66  tb=0.41
xunit15-16  15  16  unitrc1  ra=882.07  tb=0.44
xunit15-17  15  17  unitrc1  ra=3288.40  tb=0.07
xunit15-20  15  20  unitrc1  ra=2754.05  tb=0.12
xunit15-23  15  23  unitrc1  ra=1878.78  tb=0.38
xunit15-24  15  24  unitrc1  ra=3377.27  tb=0.17
xunit15-27  15  27  unitrc1  ra=6012.34  tb=0.06
xunit15-33  15  33  unitrc1  ra=3940.91  tb=0.10
xunit15-34  15  34  unitrc1  ra=9910.35  tb=0.36
xunit15-36  15  36  unitrc1  ra=1337.73  tb=0.05
xunit15-39  15  39  unitrc1  ra=4331.64  tb=0.10
xunit15-40  15  40  unitrc1  ra=6272.22  tb=0.04
xunit15-41  15  41  unitrc1  ra=267.31  tb=0.37
xunit15-42  15  42  unitrc1  ra=4268.35  tb=0.27
xunit15-43  15  43  unitrc1  ra=5257.40  tb=0.21

xunit16-1  16  1  unitrc1  ra=5883.90  tb=0.22
xunit16-2  16  2  unitrc1  ra=2515.84  tb=0.48
xunit16-3  16  3  unitrc1  ra=1513.67  tb=0.15
xunit16-5  16  5  unitrc1  ra=6241.79  tb=0.20
xunit16-8  16  8  unitrc1  ra=1020.01  tb=0.36
xunit16-10  16  10  unitrc1  ra=4365.88  tb=0.01
xunit16-13  16  13  unitrc1  ra=6871.32  tb=0.31
xunit16-17  16  17  unitrc1  ra=6885.16  tb=0.43
xunit16-20  16  20  unitrc1  ra=886.23  tb=0.24
xunit16-21  16  21  unitrc1  ra=1476.25  tb=0.07
xunit16-22  16  22  unitrc1  ra=3532.07  tb=0.41
xunit16-25  16  25  unitrc1  ra=5109.35  tb=0.22
xunit16-28  16  28  unitrc1  ra=2815.97  tb=0.09
xunit16-29  16  29  unitrc1  ra=5895.97  tb=0.37
xunit16-30  16  30  unitrc1  ra=7321.60  tb=0.07
xunit16-31  16  31  unitrc1  ra=7084.00  tb=0.47
xunit16-32  16  32  unitrc1  ra=878.66  tb=0.36
xunit16-34  16  34  unitrc1  ra=1810.25  tb=0.34
xunit16-35  16  35  unitrc1  ra=6248.37  tb=0.14
xunit16-36  16  36  unitrc1  ra=8946.22  tb=0.05
xunit16-37  16  37  unitrc1  ra=6650.19  tb=0.21
xunit16-39  16  39  unitrc1  ra=5736.65  tb=0.36
xunit16-40  16  40  unitrc1  ra=6139.41  tb=0.15
xunit16-44  16  44  unitrc1  ra=3789.13  tb=0.32
xunit16-45  16  45  unitrc1  ra=5439.45  tb=0.22
xunit16-47  16  47  unitrc1  ra=893.32  tb=0.16
xunit16-48  16  48  unitrc1  ra=864.71  tb=0.16
xunit16-49  16  49  unitrc1  ra=4118.46  tb=0.30
xunit16-50  16  50  unitrc1  ra=6382.20  tb=0.36

xunit17-5  17  5  unitrc1  ra=2717.00  tb=0.12
xunit17-6  17  6  unitrc1  ra=3687.47  tb=0.41
xunit17-7  17  7  unitrc1  ra=5495.88  tb=0.10
xunit17-8  17  8  unitrc1  ra=1783.85  tb=0.19
xunit17-12  17  12  unitrc1  ra=2194.90  tb=0.06
xunit17-13  17  13  unitrc1  ra=2163.70  tb=0.43
xunit17-14  17  14  unitrc1  ra=6354.28  tb=0.41
xunit17-15  17  15  unitrc1  ra=1175.75  tb=0.20
xunit17-18  17  18  unitrc1  ra=259.80  tb=0.45
xunit17-22  17  22  unitrc1  ra=8705.16  tb=0.38
xunit17-23  17  23  unitrc1  ra=5508.29  tb=0.14
xunit17-28  17  28  unitrc1  ra=3132.68  tb=0.28
xunit17-33  17  33  unitrc1  ra=1606.86  tb=0.39
xunit17-34  17  34  unitrc1  ra=9402.96  tb=0.48
xunit17-35  17  35  unitrc1  ra=8851.88  tb=0.20
xunit17-39  17  39  unitrc1  ra=4942.91  tb=0.36
xunit17-40  17  40  unitrc1  ra=1766.95  tb=0.27
xunit17-42  17  42  unitrc1  ra=5344.00  tb=0.06
xunit17-43  17  43  unitrc1  ra=8158.36  tb=0.34
xunit17-44  17  44  unitrc1  ra=701.62  tb=0.44
xunit17-45  17  45  unitrc1  ra=3108.74  tb=0.33
xunit17-46  17  46  unitrc1  ra=668.18  tb=0.17
xunit17-50  17  50  unitrc1  ra=1015.09  tb=0.32

xunit18-1  18  1  unitrc1  ra=2658.14  tb=0.28
xunit18-2  18  2  unitrc1  ra=7422.93  tb=0.29
xunit18-3  18  3  unitrc1  ra=8266.98  tb=0.42
xunit18-4  18  4  unitrc1  ra=808.97  tb=0.47
xunit18-5  18  5  unitrc1  ra=1624.76  tb=0.39
xunit18-6  18  6  unitrc1  ra=2285.18  tb=0.11
xunit18-7  18  7  unitrc1  ra=5657.36  tb=0.36
xunit18-9  18  9  unitrc1  ra=557.08  tb=0.12
xunit18-12  18  12  unitrc1  ra=1943.70  tb=0.20
xunit18-13  18  13  unitrc1  ra=5661.83  tb=0.16
xunit18-15  18  15  unitrc1  ra=1907.20  tb=0.15
xunit18-17  18  17  unitrc1  ra=6940.16  tb=0.36
xunit18-18  18  18  unitrc1  ra=4529.99  tb=0.10
xunit18-19  18  19  unitrc1  ra=5904.93  tb=0.10
xunit18-20  18  20  unitrc1  ra=7673.02  tb=0.21
xunit18-22  18  22  unitrc1  ra=2776.59  tb=0.02
xunit18-26  18  26  unitrc1  ra=2398.21  tb=0.13
xunit18-27  18  27  unitrc1  ra=7375.32  tb=0.39
xunit18-28  18  28  unitrc1  ra=1796.50  tb=0.45
xunit18-29  18  29  unitrc1  ra=2088.86  tb=0.26
xunit18-30  18  30  unitrc1  ra=1157.82  tb=0.20
xunit18-32  18  32  unitrc1  ra=6622.81  tb=0.48
xunit18-34  18  34  unitrc1  ra=964.16  tb=0.25
xunit18-35  18  35  unitrc1  ra=2925.07  tb=0.43
xunit18-38  18  38  unitrc1  ra=3405.27  tb=0.06
xunit18-40  18  40  unitrc1  ra=9914.81  tb=0.08
xunit18-41  18  41  unitrc1  ra=5789.03  tb=0.08
xunit18-42  18  42  unitrc1  ra=5290.52  tb=0.42
xunit18-44  18  44  unitrc1  ra=3770.62  tb=0.22
xunit18-45  18  45  unitrc1  ra=5318.79  tb=0.32

xunit19-1  19  1  unitrc1  ra=1498.05  tb=0.00
xunit19-4  19  4  unitrc1  ra=2000.51  tb=0.46
xunit19-5  19  5  unitrc1  ra=6006.72  tb=0.09
xunit19-7  19  7  unitrc1  ra=5787.82  tb=0.08
xunit19-8  19  8  unitrc1  ra=4565.41  tb=0.16
xunit19-13  19  13  unitrc1  ra=1860.78  tb=0.17
xunit19-14  19  14  unitrc1  ra=3245.87  tb=0.31
xunit19-15  19  15  unitrc1  ra=5018.14  tb=0.40
xunit19-16  19  16  unitrc1  ra=3524.44  tb=0.24
xunit19-17  19  17  unitrc1  ra=8660.19  tb=0.19
xunit19-20  19  20  unitrc1  ra=2879.55  tb=0.11
xunit19-22  19  22  unitrc1  ra=4406.85  tb=0.45
xunit19-23  19  23  unitrc1  ra=3190.08  tb=0.10
xunit19-24  19  24  unitrc1  ra=4849.17  tb=0.47
xunit19-25  19  25  unitrc1  ra=1294.79  tb=0.26
xunit19-26  19  26  unitrc1  ra=462.86  tb=0.16
xunit19-27  19  27  unitrc1  ra=7878.21  tb=0.09
xunit19-28  19  28  unitrc1  ra=8909.80  tb=0.10
xunit19-29  19  29  unitrc1  ra=6474.51  tb=0.36
xunit19-30  19  30  unitrc1  ra=3269.55  tb=0.15
xunit19-31  19  31  unitrc1  ra=4816.15  tb=0.17
xunit19-33  19  33  unitrc1  ra=2766.87  tb=0.28
xunit19-36  19  36  unitrc1  ra=142.99  tb=0.20
xunit19-37  19  37  unitrc1  ra=251.93  tb=0.11
xunit19-39  19  39  unitrc1  ra=5531.45  tb=0.30
xunit19-44  19  44  unitrc1  ra=1070.09  tb=0.17
xunit19-48  19  48  unitrc1  ra=7093.80  tb=0.20
xunit19-50  19  50  unitrc1  ra=8174.29  tb=0.18

xunit20-1  20  1  unitrc1  ra=1938.45  tb=0.29
xunit20-4  20  4  unitrc1  ra=2679.41  tb=0.19
xunit20-8  20  8  unitrc1  ra=170.29  tb=0.36
xunit20-9  20  9  unitrc1  ra=9075.90  tb=0.49
xunit20-13  20  13  unitrc1  ra=3130.54  tb=0.02
xunit20-15  20  15  unitrc1  ra=4894.66  tb=0.11
xunit20-17  20  17  unitrc1  ra=9610.26  tb=0.17
xunit20-18  20  18  unitrc1  ra=4037.78  tb=0.27
xunit20-19  20  19  unitrc1  ra=1377.38  tb=0.14
xunit20-20  20  20  unitrc1  ra=8462.03  tb=0.36
xunit20-21  20  21  unitrc1  ra=1267.84  tb=0.10
xunit20-22  20  22  unitrc1  ra=734.30  tb=0.16
xunit20-23  20  23  unitrc1  ra=1585.32  tb=0.01
xunit20-24  20  24  unitrc1  ra=6732.11  tb=0.34
xunit20-25  20  25  unitrc1  ra=1620.39  tb=0.16
xunit20-26  20  26  unitrc1  ra=9480.90  tb=0.43
xunit20-28  20  28  unitrc1  ra=1075.40  tb=0.16
xunit20-32  20  32  unitrc1  ra=2393.85  tb=0.19
xunit20-33  20  33  unitrc1  ra=3419.70  tb=0.43
xunit20-34  20  34  unitrc1  ra=6436.57  tb=0.40
xunit20-35  20  35  unitrc1  ra=6649.46  tb=0.46
xunit20-38  20  38  unitrc1  ra=4846.97  tb=0.50
xunit20-40  20  40  unitrc1  ra=5338.29  tb=0.25
xunit20-43  20  43  unitrc1  ra=3815.50  tb=0.41
xunit20-44  20  44  unitrc1  ra=4623.01  tb=0.09
xunit20-45  20  45  unitrc1  ra=2410.61  tb=0.11
xunit20-46  20  46  unitrc1  ra=8583.31  tb=0.42
xunit20-48  20  48  unitrc1  ra=1435.17  tb=0.17
xunit20-49  20  49  unitrc1  ra=3565.32  tb=0.08
xunit20-50  20  50  unitrc1  ra=2809.26  tb=0.27

xunit21-2  21  2  unitrc1  ra=3141.85  tb=0.41
xunit21-7  21  7  unitrc1  ra=3613.51  tb=0.38
xunit21-10  21  10  unitrc1  ra=7967.16  tb=0.04
xunit21-13  21  13  unitrc1  ra=3346.67  tb=0.47
xunit21-14  21  14  unitrc1  ra=2346.04  tb=0.38
xunit21-16  21  16  unitrc1  ra=122.81  tb=0.40
xunit21-17  21  17  unitrc1  ra=9330.75  tb=0.47
xunit21-18  21  18  unitrc1  ra=2771.92  tb=0.22
xunit21-19  21  19  unitrc1  ra=5662.95  tb=0.28
xunit21-22  21  22  unitrc1  ra=3238.16  tb=0.11
xunit21-23  21  23  unitrc1  ra=4078.50  tb=0.30
xunit21-24  21  24  unitrc1  ra=2699.41  tb=0.18
xunit21-25  21  25  unitrc1  ra=780.61  tb=0.34
xunit21-26  21  26  unitrc1  ra=1956.65  tb=0.24
xunit21-29  21  29  unitrc1  ra=810.97  tb=0.26
xunit21-30  21  30  unitrc1  ra=5266.92  tb=0.20
xunit21-31  21  31  unitrc1  ra=3392.68  tb=0.23
xunit21-33  21  33  unitrc1  ra=1935.58  tb=0.03
xunit21-35  21  35  unitrc1  ra=1712.35  tb=0.29
xunit21-36  21  36  unitrc1  ra=3254.50  tb=0.10
xunit21-37  21  37  unitrc1  ra=5411.89  tb=0.39
xunit21-38  21  38  unitrc1  ra=8338.33  tb=0.46
xunit21-39  21  39  unitrc1  ra=7439.46  tb=0.13
xunit21-41  21  41  unitrc1  ra=1011.62  tb=0.49
xunit21-42  21  42  unitrc1  ra=2546.53  tb=0.25
xunit21-47  21  47  unitrc1  ra=7790.80  tb=0.41
xunit21-48  21  48  unitrc1  ra=1160.96  tb=0.18
xunit21-49  21  49  unitrc1  ra=2587.41  tb=0.44

xunit22-1  22  1  unitrc1  ra=8947.57  tb=0.39
xunit22-2  22  2  unitrc1  ra=6718.61  tb=0.45
xunit22-3  22  3  unitrc1  ra=5688.64  tb=0.39
xunit22-5  22  5  unitrc1  ra=6300.29  tb=0.34
xunit22-7  22  7  unitrc1  ra=6445.57  tb=0.01
xunit22-8  22  8  unitrc1  ra=5331.27  tb=0.43
xunit22-9  22  9  unitrc1  ra=9806.66  tb=0.36
xunit22-14  22  14  unitrc1  ra=4813.26  tb=0.34
xunit22-15  22  15  unitrc1  ra=7392.02  tb=0.24
xunit22-16  22  16  unitrc1  ra=1987.60  tb=0.45
xunit22-18  22  18  unitrc1  ra=6470.33  tb=0.04
xunit22-20  22  20  unitrc1  ra=6353.72  tb=0.13
xunit22-23  22  23  unitrc1  ra=3232.17  tb=0.27
xunit22-25  22  25  unitrc1  ra=8211.76  tb=0.32
xunit22-31  22  31  unitrc1  ra=6317.00  tb=0.31
xunit22-33  22  33  unitrc1  ra=9644.94  tb=0.27
xunit22-35  22  35  unitrc1  ra=3155.23  tb=0.30
xunit22-37  22  37  unitrc1  ra=7780.95  tb=0.28
xunit22-38  22  38  unitrc1  ra=3209.76  tb=0.24
xunit22-39  22  39  unitrc1  ra=832.45  tb=0.02
xunit22-40  22  40  unitrc1  ra=2824.59  tb=0.05
xunit22-41  22  41  unitrc1  ra=3739.34  tb=0.31
xunit22-42  22  42  unitrc1  ra=7481.23  tb=0.45
xunit22-43  22  43  unitrc1  ra=3824.79  tb=0.32
xunit22-44  22  44  unitrc1  ra=6163.52  tb=0.25
xunit22-47  22  47  unitrc1  ra=4847.40  tb=0.31
xunit22-48  22  48  unitrc1  ra=3402.77  tb=0.01
xunit22-49  22  49  unitrc1  ra=4636.64  tb=0.27

xunit23-1  23  1  unitrc1  ra=382.21  tb=0.24
xunit23-2  23  2  unitrc1  ra=6817.02  tb=0.11
xunit23-5  23  5  unitrc1  ra=3212.99  tb=0.41
xunit23-8  23  8  unitrc1  ra=4279.32  tb=0.36
xunit23-9  23  9  unitrc1  ra=2648.83  tb=0.16
xunit23-10  23  10  unitrc1  ra=9769.56  tb=0.42
xunit23-11  23  11  unitrc1  ra=4050.75  tb=0.26
xunit23-12  23  12  unitrc1  ra=4044.84  tb=0.47
xunit23-13  23  13  unitrc1  ra=7921.16  tb=0.40
xunit23-17  23  17  unitrc1  ra=6571.60  tb=0.32
xunit23-19  23  19  unitrc1  ra=110.94  tb=0.19
xunit23-20  23  20  unitrc1  ra=6876.23  tb=0.36
xunit23-21  23  21  unitrc1  ra=8653.35  tb=0.28
xunit23-22  23  22  unitrc1  ra=8378.19  tb=0.40
xunit23-24  23  24  unitrc1  ra=9805.55  tb=0.26
xunit23-25  23  25  unitrc1  ra=3457.16  tb=0.43
xunit23-26  23  26  unitrc1  ra=5160.13  tb=0.26
xunit23-27  23  27  unitrc1  ra=4462.70  tb=0.09
xunit23-28  23  28  unitrc1  ra=1949.32  tb=0.28
xunit23-29  23  29  unitrc1  ra=5174.84  tb=0.09
xunit23-31  23  31  unitrc1  ra=4997.96  tb=0.29
xunit23-35  23  35  unitrc1  ra=3527.05  tb=0.22
xunit23-37  23  37  unitrc1  ra=1508.97  tb=0.40
xunit23-38  23  38  unitrc1  ra=5409.66  tb=0.03
xunit23-39  23  39  unitrc1  ra=4340.48  tb=0.34
xunit23-40  23  40  unitrc1  ra=1581.50  tb=0.49
xunit23-41  23  41  unitrc1  ra=395.79  tb=0.33
xunit23-44  23  44  unitrc1  ra=3182.38  tb=0.20
xunit23-47  23  47  unitrc1  ra=3966.51  tb=0.34
xunit23-50  23  50  unitrc1  ra=6729.38  tb=0.44

xunit24-1  24  1  unitrc1  ra=5421.15  tb=0.02
xunit24-4  24  4  unitrc1  ra=2990.28  tb=0.03
xunit24-5  24  5  unitrc1  ra=1444.38  tb=0.13
xunit24-7  24  7  unitrc1  ra=5301.47  tb=0.18
xunit24-8  24  8  unitrc1  ra=1399.91  tb=0.16
xunit24-9  24  9  unitrc1  ra=5985.78  tb=0.25
xunit24-11  24  11  unitrc1  ra=9389.19  tb=0.33
xunit24-13  24  13  unitrc1  ra=3052.41  tb=0.16
xunit24-14  24  14  unitrc1  ra=322.46  tb=0.45
xunit24-15  24  15  unitrc1  ra=2925.14  tb=0.23
xunit24-16  24  16  unitrc1  ra=1593.81  tb=0.44
xunit24-17  24  17  unitrc1  ra=6653.26  tb=0.11
xunit24-18  24  18  unitrc1  ra=3375.06  tb=0.01
xunit24-19  24  19  unitrc1  ra=809.22  tb=0.12
xunit24-20  24  20  unitrc1  ra=3124.96  tb=0.23
xunit24-21  24  21  unitrc1  ra=4945.34  tb=0.18
xunit24-22  24  22  unitrc1  ra=7269.42  tb=0.10
xunit24-23  24  23  unitrc1  ra=2013.66  tb=0.14
xunit24-24  24  24  unitrc1  ra=8232.87  tb=0.26
xunit24-25  24  25  unitrc1  ra=3954.41  tb=0.31
xunit24-27  24  27  unitrc1  ra=8913.61  tb=0.16
xunit24-29  24  29  unitrc1  ra=5853.09  tb=0.43
xunit24-31  24  31  unitrc1  ra=2538.36  tb=0.22
xunit24-32  24  32  unitrc1  ra=4866.17  tb=0.13
xunit24-34  24  34  unitrc1  ra=2720.70  tb=0.15
xunit24-35  24  35  unitrc1  ra=4513.88  tb=0.21
xunit24-36  24  36  unitrc1  ra=557.32  tb=0.16
xunit24-37  24  37  unitrc1  ra=8398.31  tb=0.36
xunit24-38  24  38  unitrc1  ra=1816.80  tb=0.42
xunit24-42  24  42  unitrc1  ra=7865.96  tb=0.38
xunit24-45  24  45  unitrc1  ra=143.47  tb=0.06
xunit24-46  24  46  unitrc1  ra=2783.08  tb=0.06
xunit24-48  24  48  unitrc1  ra=4878.87  tb=0.42
xunit24-50  24  50  unitrc1  ra=2178.76  tb=0.02

xunit25-2  25  2  unitrc1  ra=1918.69  tb=0.09
xunit25-4  25  4  unitrc1  ra=3324.12  tb=0.49
xunit25-6  25  6  unitrc1  ra=5884.95  tb=0.29
xunit25-8  25  8  unitrc1  ra=9667.45  tb=0.23
xunit25-10  25  10  unitrc1  ra=2781.23  tb=0.41
xunit25-11  25  11  unitrc1  ra=3895.30  tb=0.33
xunit25-12  25  12  unitrc1  ra=6350.29  tb=0.14
xunit25-15  25  15  unitrc1  ra=2913.52  tb=0.23
xunit25-18  25  18  unitrc1  ra=5594.07  tb=0.25
xunit25-20  25  20  unitrc1  ra=6405.27  tb=0.23
xunit25-21  25  21  unitrc1  ra=5944.29  tb=0.02
xunit25-23  25  23  unitrc1  ra=5921.01  tb=0.12
xunit25-24  25  24  unitrc1  ra=3716.32  tb=0.38
xunit25-25  25  25  unitrc1  ra=9226.72  tb=0.15
xunit25-26  25  26  unitrc1  ra=5241.25  tb=0.24
xunit25-28  25  28  unitrc1  ra=596.90  tb=0.23
xunit25-30  25  30  unitrc1  ra=1630.04  tb=0.09
xunit25-31  25  31  unitrc1  ra=4522.25  tb=0.21
xunit25-34  25  34  unitrc1  ra=4020.31  tb=0.05
xunit25-35  25  35  unitrc1  ra=4957.83  tb=0.35
xunit25-36  25  36  unitrc1  ra=669.86  tb=0.47
xunit25-39  25  39  unitrc1  ra=2407.37  tb=0.17
xunit25-40  25  40  unitrc1  ra=5315.34  tb=0.23
xunit25-41  25  41  unitrc1  ra=2967.97  tb=0.17
xunit25-44  25  44  unitrc1  ra=6019.91  tb=0.36
xunit25-46  25  46  unitrc1  ra=5767.24  tb=0.28
xunit25-47  25  47  unitrc1  ra=4534.52  tb=0.47

xunit26-2  26  2  unitrc1  ra=6476.79  tb=0.32
xunit26-4  26  4  unitrc1  ra=748.16  tb=0.33
xunit26-5  26  5  unitrc1  ra=4880.98  tb=0.27
xunit26-6  26  6  unitrc1  ra=6123.50  tb=0.33
xunit26-9  26  9  unitrc1  ra=2625.83  tb=0.24
xunit26-16  26  16  unitrc1  ra=2665.06  tb=0.18
xunit26-17  26  17  unitrc1  ra=5739.41  tb=0.38
xunit26-21  26  21  unitrc1  ra=6351.28  tb=0.20
xunit26-24  26  24  unitrc1  ra=9915.19  tb=0.41
xunit26-25  26  25  unitrc1  ra=845.16  tb=0.20
xunit26-26  26  26  unitrc1  ra=1365.41  tb=0.13
xunit26-27  26  27  unitrc1  ra=7361.75  tb=0.05
xunit26-29  26  29  unitrc1  ra=5628.09  tb=0.21
xunit26-30  26  30  unitrc1  ra=9321.99  tb=0.11
xunit26-31  26  31  unitrc1  ra=5132.84  tb=0.32
xunit26-32  26  32  unitrc1  ra=4693.92  tb=0.24
xunit26-34  26  34  unitrc1  ra=2659.54  tb=0.07
xunit26-35  26  35  unitrc1  ra=3394.27  tb=0.08
xunit26-36  26  36  unitrc1  ra=3624.51  tb=0.19
xunit26-37  26  37  unitrc1  ra=4907.74  tb=0.30
xunit26-38  26  38  unitrc1  ra=4516.85  tb=0.10
xunit26-39  26  39  unitrc1  ra=2592.01  tb=0.06
xunit26-40  26  40  unitrc1  ra=1492.68  tb=0.34
xunit26-41  26  41  unitrc1  ra=2859.55  tb=0.36
xunit26-43  26  43  unitrc1  ra=1184.21  tb=0.40
xunit26-44  26  44  unitrc1  ra=6120.62  tb=0.04
xunit26-45  26  45  unitrc1  ra=5017.29  tb=0.49
xunit26-47  26  47  unitrc1  ra=5697.92  tb=0.10
xunit26-48  26  48  unitrc1  ra=2503.40  tb=0.34
xunit26-50  26  50  unitrc1  ra=2438.71  tb=0.09

xunit27-2  27  2  unitrc1  ra=1621.04  tb=0.33
xunit27-6  27  6  unitrc1  ra=6175.52  tb=0.12
xunit27-7  27  7  unitrc1  ra=8672.25  tb=0.20
xunit27-8  27  8  unitrc1  ra=7687.00  tb=0.44
xunit27-9  27  9  unitrc1  ra=2837.56  tb=0.09
xunit27-10  27  10  unitrc1  ra=582.75  tb=0.28
xunit27-11  27  11  unitrc1  ra=538.48  tb=0.33
xunit27-13  27  13  unitrc1  ra=6217.63  tb=0.23
xunit27-16  27  16  unitrc1  ra=8189.50  tb=0.14
xunit27-17  27  17  unitrc1  ra=6404.82  tb=0.23
xunit27-19  27  19  unitrc1  ra=3190.62  tb=0.07
xunit27-20  27  20  unitrc1  ra=2022.05  tb=0.27
xunit27-21  27  21  unitrc1  ra=3610.94  tb=0.25
xunit27-22  27  22  unitrc1  ra=4496.67  tb=0.02
xunit27-24  27  24  unitrc1  ra=8312.70  tb=0.40
xunit27-25  27  25  unitrc1  ra=4891.36  tb=0.04
xunit27-26  27  26  unitrc1  ra=4703.17  tb=0.20
xunit27-27  27  27  unitrc1  ra=6931.74  tb=0.09
xunit27-28  27  28  unitrc1  ra=7129.37  tb=0.01
xunit27-29  27  29  unitrc1  ra=1152.68  tb=0.15
xunit27-31  27  31  unitrc1  ra=5141.70  tb=0.15
xunit27-32  27  32  unitrc1  ra=8811.90  tb=0.10
xunit27-33  27  33  unitrc1  ra=2159.67  tb=0.15
xunit27-34  27  34  unitrc1  ra=1307.79  tb=0.39
xunit27-36  27  36  unitrc1  ra=1656.49  tb=0.24
xunit27-37  27  37  unitrc1  ra=4302.78  tb=0.17
xunit27-39  27  39  unitrc1  ra=4878.09  tb=0.34
xunit27-40  27  40  unitrc1  ra=3570.88  tb=0.09
xunit27-42  27  42  unitrc1  ra=3630.76  tb=0.44
xunit27-43  27  43  unitrc1  ra=248.73  tb=0.12
xunit27-44  27  44  unitrc1  ra=8410.49  tb=0.11
xunit27-45  27  45  unitrc1  ra=7523.50  tb=0.08
xunit27-46  27  46  unitrc1  ra=2658.57  tb=0.35

xunit28-1  28  1  unitrc1  ra=8436.36  tb=0.27
xunit28-4  28  4  unitrc1  ra=5010.91  tb=0.24
xunit28-6  28  6  unitrc1  ra=2691.07  tb=0.31
xunit28-11  28  11  unitrc1  ra=9651.48  tb=0.50
xunit28-12  28  12  unitrc1  ra=827.93  tb=0.29
xunit28-14  28  14  unitrc1  ra=6992.72  tb=0.20
xunit28-17  28  17  unitrc1  ra=4974.64  tb=0.49
xunit28-22  28  22  unitrc1  ra=6669.80  tb=0.26
xunit28-24  28  24  unitrc1  ra=9604.92  tb=0.36
xunit28-28  28  28  unitrc1  ra=5004.60  tb=0.49
xunit28-29  28  29  unitrc1  ra=6534.21  tb=0.34
xunit28-30  28  30  unitrc1  ra=3666.85  tb=0.07
xunit28-31  28  31  unitrc1  ra=6323.42  tb=0.14
xunit28-32  28  32  unitrc1  ra=5275.69  tb=0.18
xunit28-36  28  36  unitrc1  ra=1159.69  tb=0.32
xunit28-37  28  37  unitrc1  ra=2577.62  tb=0.01
xunit28-39  28  39  unitrc1  ra=3164.23  tb=0.35
xunit28-41  28  41  unitrc1  ra=6269.71  tb=0.01
xunit28-42  28  42  unitrc1  ra=3692.82  tb=0.35
xunit28-43  28  43  unitrc1  ra=831.63  tb=0.09
xunit28-45  28  45  unitrc1  ra=2831.59  tb=0.44
xunit28-46  28  46  unitrc1  ra=4523.05  tb=0.16
xunit28-47  28  47  unitrc1  ra=5154.36  tb=0.45
xunit28-48  28  48  unitrc1  ra=9890.94  tb=0.26
xunit28-50  28  50  unitrc1  ra=702.70  tb=0.38

xunit29-1  29  1  unitrc1  ra=6182.01  tb=0.46
xunit29-2  29  2  unitrc1  ra=1764.22  tb=0.24
xunit29-9  29  9  unitrc1  ra=1795.15  tb=0.24
xunit29-12  29  12  unitrc1  ra=3266.75  tb=0.26
xunit29-13  29  13  unitrc1  ra=721.14  tb=0.14
xunit29-15  29  15  unitrc1  ra=4943.40  tb=0.27
xunit29-16  29  16  unitrc1  ra=1269.35  tb=0.24
xunit29-17  29  17  unitrc1  ra=2578.21  tb=0.01
xunit29-18  29  18  unitrc1  ra=5982.01  tb=0.21
xunit29-21  29  21  unitrc1  ra=4071.44  tb=0.47
xunit29-22  29  22  unitrc1  ra=4247.92  tb=0.11
xunit29-26  29  26  unitrc1  ra=1734.03  tb=0.36
xunit29-27  29  27  unitrc1  ra=9827.26  tb=0.16
xunit29-30  29  30  unitrc1  ra=4529.46  tb=0.47
xunit29-32  29  32  unitrc1  ra=4767.67  tb=0.29
xunit29-34  29  34  unitrc1  ra=8486.41  tb=0.15
xunit29-35  29  35  unitrc1  ra=3103.00  tb=0.29
xunit29-37  29  37  unitrc1  ra=213.28  tb=0.38
xunit29-38  29  38  unitrc1  ra=5022.09  tb=0.26
xunit29-39  29  39  unitrc1  ra=4248.96  tb=0.18
xunit29-41  29  41  unitrc1  ra=2192.58  tb=0.47
xunit29-42  29  42  unitrc1  ra=2518.78  tb=0.20
xunit29-45  29  45  unitrc1  ra=8100.72  tb=0.07
xunit29-47  29  47  unitrc1  ra=279.58  tb=0.09

xunit30-2  30  2  unitrc1  ra=2461.98  tb=0.18
xunit30-3  30  3  unitrc1  ra=5209.91  tb=0.18
xunit30-5  30  5  unitrc1  ra=996.77  tb=0.25
xunit30-6  30  6  unitrc1  ra=723.32  tb=0.21
xunit30-8  30  8  unitrc1  ra=8489.76  tb=0.45
xunit30-9  30  9  unitrc1  ra=1306.62  tb=0.28
xunit30-10  30  10  unitrc1  ra=4475.92  tb=0.01
xunit30-12  30  12  unitrc1  ra=6685.06  tb=0.42
xunit30-13  30  13  unitrc1  ra=5514.39  tb=0.34
xunit30-16  30  16  unitrc1  ra=4832.89  tb=0.05
xunit30-17  30  17  unitrc1  ra=3914.32  tb=0.14
xunit30-20  30  20  unitrc1  ra=1325.59  tb=0.03
xunit30-21  30  21  unitrc1  ra=4155.96  tb=0.35
xunit30-22  30  22  unitrc1  ra=6823.54  tb=0.35
xunit30-23  30  23  unitrc1  ra=9118.57  tb=0.22
xunit30-24  30  24  unitrc1  ra=1742.54  tb=0.02
xunit30-25  30  25  unitrc1  ra=121.60  tb=0.36
xunit30-26  30  26  unitrc1  ra=3900.65  tb=0.29
xunit30-27  30  27  unitrc1  ra=4124.74  tb=0.43
xunit30-28  30  28  unitrc1  ra=3263.86  tb=0.20
xunit30-31  30  31  unitrc1  ra=7663.91  tb=0.47
xunit30-34  30  34  unitrc1  ra=3736.79  tb=0.37
xunit30-37  30  37  unitrc1  ra=217.65  tb=0.31
xunit30-38  30  38  unitrc1  ra=8699.53  tb=0.06
xunit30-39  30  39  unitrc1  ra=6815.86  tb=0.31
xunit30-40  30  40  unitrc1  ra=1906.35  tb=0.37
xunit30-42  30  42  unitrc1  ra=5613.87  tb=0.36
xunit30-43  30  43  unitrc1  ra=895.21  tb=0.44
xunit30-45  30  45  unitrc1  ra=5453.59  tb=0.50
xunit30-46  30  46  unitrc1  ra=6304.88  tb=0.32
xunit30-47  30  47  unitrc1  ra=3832.19  tb=0.27
xunit30-49  30  49  unitrc1  ra=9693.01  tb=0.06
xunit30-50  30  50  unitrc1  ra=2988.50  tb=0.27

xunit31-1  31  1  unitrc1  ra=3206.19  tb=0.29
xunit31-4  31  4  unitrc1  ra=3463.45  tb=0.17
xunit31-8  31  8  unitrc1  ra=1189.69  tb=0.30
xunit31-9  31  9  unitrc1  ra=4608.43  tb=0.36
xunit31-10  31  10  unitrc1  ra=5855.36  tb=0.04
xunit31-11  31  11  unitrc1  ra=5760.30  tb=0.17
xunit31-12  31  12  unitrc1  ra=6420.35  tb=0.23
xunit31-13  31  13  unitrc1  ra=1709.15  tb=0.12
xunit31-16  31  16  unitrc1  ra=851.71  tb=0.35
xunit31-18  31  18  unitrc1  ra=8766.05  tb=0.31
xunit31-21  31  21  unitrc1  ra=2705.95  tb=0.26
xunit31-22  31  22  unitrc1  ra=2063.50  tb=0.12
xunit31-23  31  23  unitrc1  ra=5724.71  tb=0.20
xunit31-25  31  25  unitrc1  ra=9667.72  tb=0.45
xunit31-26  31  26  unitrc1  ra=6228.12  tb=0.15
xunit31-30  31  30  unitrc1  ra=6362.77  tb=0.23
xunit31-32  31  32  unitrc1  ra=8648.13  tb=0.07
xunit31-33  31  33  unitrc1  ra=3518.27  tb=0.40
xunit31-34  31  34  unitrc1  ra=2261.52  tb=0.05
xunit31-35  31  35  unitrc1  ra=6219.32  tb=0.44
xunit31-36  31  36  unitrc1  ra=6055.79  tb=0.25
xunit31-38  31  38  unitrc1  ra=8476.51  tb=0.49
xunit31-40  31  40  unitrc1  ra=1952.12  tb=0.42
xunit31-41  31  41  unitrc1  ra=420.55  tb=0.09
xunit31-42  31  42  unitrc1  ra=2126.97  tb=0.21
xunit31-44  31  44  unitrc1  ra=4488.72  tb=0.41
xunit31-45  31  45  unitrc1  ra=4788.98  tb=0.24
xunit31-46  31  46  unitrc1  ra=2128.57  tb=0.36
xunit31-47  31  47  unitrc1  ra=4962.31  tb=0.14
xunit31-48  31  48  unitrc1  ra=8861.53  tb=0.42
xunit31-49  31  49  unitrc1  ra=3629.57  tb=0.20

xunit32-2  32  2  unitrc1  ra=6204.13  tb=0.40
xunit32-5  32  5  unitrc1  ra=4617.14  tb=0.37
xunit32-6  32  6  unitrc1  ra=358.86  tb=0.26
xunit32-7  32  7  unitrc1  ra=2553.02  tb=0.17
xunit32-8  32  8  unitrc1  ra=6606.52  tb=0.28
xunit32-10  32  10  unitrc1  ra=6203.64  tb=0.25
xunit32-11  32  11  unitrc1  ra=723.87  tb=0.25
xunit32-12  32  12  unitrc1  ra=3281.77  tb=0.08
xunit32-13  32  13  unitrc1  ra=3541.08  tb=0.35
xunit32-14  32  14  unitrc1  ra=758.43  tb=0.26
xunit32-15  32  15  unitrc1  ra=1222.72  tb=0.14
xunit32-16  32  16  unitrc1  ra=8121.70  tb=0.16
xunit32-21  32  21  unitrc1  ra=6314.26  tb=0.44
xunit32-24  32  24  unitrc1  ra=1784.41  tb=0.33
xunit32-25  32  25  unitrc1  ra=5689.24  tb=0.29
xunit32-28  32  28  unitrc1  ra=5682.68  tb=0.38
xunit32-29  32  29  unitrc1  ra=3668.55  tb=0.15
xunit32-30  32  30  unitrc1  ra=1314.53  tb=0.08
xunit32-31  32  31  unitrc1  ra=4173.91  tb=0.05
xunit32-33  32  33  unitrc1  ra=7949.05  tb=0.08
xunit32-34  32  34  unitrc1  ra=2569.57  tb=0.18
xunit32-36  32  36  unitrc1  ra=722.42  tb=0.30
xunit32-38  32  38  unitrc1  ra=4333.21  tb=0.41
xunit32-39  32  39  unitrc1  ra=3453.30  tb=0.28
xunit32-43  32  43  unitrc1  ra=1770.90  tb=0.23
xunit32-46  32  46  unitrc1  ra=8180.84  tb=0.20
xunit32-48  32  48  unitrc1  ra=2619.41  tb=0.08
xunit32-49  32  49  unitrc1  ra=8454.80  tb=0.40
xunit32-50  32  50  unitrc1  ra=4460.71  tb=0.40

xunit33-1  33  1  unitrc1  ra=1096.00  tb=0.24
xunit33-3  33  3  unitrc1  ra=5524.01  tb=0.26
xunit33-4  33  4  unitrc1  ra=2150.61  tb=0.38
xunit33-5  33  5  unitrc1  ra=4422.52  tb=0.35
xunit33-8  33  8  unitrc1  ra=6181.07  tb=0.37
xunit33-10  33  10  unitrc1  ra=2737.08  tb=0.26
xunit33-11  33  11  unitrc1  ra=156.52  tb=0.32
xunit33-12  33  12  unitrc1  ra=5894.26  tb=0.46
xunit33-13  33  13  unitrc1  ra=1251.19  tb=0.36
xunit33-14  33  14  unitrc1  ra=6041.84  tb=0.11
xunit33-15  33  15  unitrc1  ra=137.95  tb=0.04
xunit33-16  33  16  unitrc1  ra=3393.74  tb=0.38
xunit33-17  33  17  unitrc1  ra=6928.95  tb=0.02
xunit33-19  33  19  unitrc1  ra=3728.91  tb=0.39
xunit33-21  33  21  unitrc1  ra=447.93  tb=0.44
xunit33-22  33  22  unitrc1  ra=4347.47  tb=0.24
xunit33-23  33  23  unitrc1  ra=5955.22  tb=0.07
xunit33-24  33  24  unitrc1  ra=2124.48  tb=0.05
xunit33-26  33  26  unitrc1  ra=4429.85  tb=0.45
xunit33-30  33  30  unitrc1  ra=2728.95  tb=0.38
xunit33-33  33  33  unitrc1  ra=1827.15  tb=0.48
xunit33-34  33  34  unitrc1  ra=4466.49  tb=0.23
xunit33-37  33  37  unitrc1  ra=3889.61  tb=0.36
xunit33-39  33  39  unitrc1  ra=1030.43  tb=0.28
xunit33-41  33  41  unitrc1  ra=3360.28  tb=0.50
xunit33-42  33  42  unitrc1  ra=6181.26  tb=0.25
xunit33-43  33  43  unitrc1  ra=3931.83  tb=0.04
xunit33-44  33  44  unitrc1  ra=543.88  tb=0.36
xunit33-45  33  45  unitrc1  ra=6636.91  tb=0.40
xunit33-46  33  46  unitrc1  ra=7313.03  tb=0.01
xunit33-47  33  47  unitrc1  ra=600.36  tb=0.44
xunit33-48  33  48  unitrc1  ra=4206.52  tb=0.32
xunit33-49  33  49  unitrc1  ra=4462.28  tb=0.11
xunit33-50  33  50  unitrc1  ra=292.89  tb=0.30

xunit34-1  34  1  unitrc1  ra=2606.76  tb=0.30
xunit34-2  34  2  unitrc1  ra=3703.16  tb=0.03
xunit34-3  34  3  unitrc1  ra=2212.66  tb=0.04
xunit34-7  34  7  unitrc1  ra=5025.19  tb=0.41
xunit34-8  34  8  unitrc1  ra=1913.11  tb=0.24
xunit34-9  34  9  unitrc1  ra=5998.14  tb=0.34
xunit34-10  34  10  unitrc1  ra=4213.63  tb=0.38
xunit34-18  34  18  unitrc1  ra=432.03  tb=0.23
xunit34-21  34  21  unitrc1  ra=6543.84  tb=0.14
xunit34-24  34  24  unitrc1  ra=2214.77  tb=0.48
xunit34-26  34  26  unitrc1  ra=7061.22  tb=0.06
xunit34-28  34  28  unitrc1  ra=2355.70  tb=0.20
xunit34-29  34  29  unitrc1  ra=646.68  tb=0.32
xunit34-31  34  31  unitrc1  ra=6430.91  tb=0.46
xunit34-32  34  32  unitrc1  ra=1107.15  tb=0.32
xunit34-34  34  34  unitrc1  ra=5411.36  tb=0.21
xunit34-35  34  35  unitrc1  ra=2714.10  tb=0.26
xunit34-39  34  39  unitrc1  ra=4851.17  tb=0.34
xunit34-40  34  40  unitrc1  ra=4521.52  tb=0.26
xunit34-41  34  41  unitrc1  ra=6073.53  tb=0.19
xunit34-44  34  44  unitrc1  ra=8872.97  tb=0.38
xunit34-45  34  45  unitrc1  ra=8986.90  tb=0.01
xunit34-47  34  47  unitrc1  ra=2623.61  tb=0.27
xunit34-48  34  48  unitrc1  ra=7765.05  tb=0.38
xunit34-50  34  50  unitrc1  ra=5873.04  tb=0.16

xunit35-1  35  1  unitrc1  ra=6020.50  tb=0.33
xunit35-2  35  2  unitrc1  ra=5723.77  tb=0.32
xunit35-4  35  4  unitrc1  ra=1889.55  tb=0.03
xunit35-8  35  8  unitrc1  ra=415.64  tb=0.10
xunit35-10  35  10  unitrc1  ra=8004.54  tb=0.36
xunit35-13  35  13  unitrc1  ra=6220.21  tb=0.07
xunit35-15  35  15  unitrc1  ra=1185.16  tb=0.05
xunit35-16  35  16  unitrc1  ra=1511.73  tb=0.27
xunit35-17  35  17  unitrc1  ra=4210.42  tb=0.42
xunit35-20  35  20  unitrc1  ra=3016.11  tb=0.46
xunit35-21  35  21  unitrc1  ra=4643.64  tb=0.05
xunit35-28  35  28  unitrc1  ra=6623.23  tb=0.36
xunit35-30  35  30  unitrc1  ra=5769.66  tb=0.24
xunit35-32  35  32  unitrc1  ra=1833.49  tb=0.36
xunit35-33  35  33  unitrc1  ra=9038.63  tb=0.13
xunit35-34  35  34  unitrc1  ra=6124.81  tb=0.21
xunit35-36  35  36  unitrc1  ra=4517.21  tb=0.06
xunit35-37  35  37  unitrc1  ra=1420.18  tb=0.19
xunit35-39  35  39  unitrc1  ra=1011.40  tb=0.20
xunit35-41  35  41  unitrc1  ra=7635.46  tb=0.12
xunit35-42  35  42  unitrc1  ra=5681.27  tb=0.34
xunit35-43  35  43  unitrc1  ra=9528.44  tb=0.16
xunit35-44  35  44  unitrc1  ra=3722.72  tb=0.03
xunit35-45  35  45  unitrc1  ra=6591.25  tb=0.30
xunit35-47  35  47  unitrc1  ra=5368.01  tb=0.20

xunit36-1  36  1  unitrc1  ra=102.52  tb=0.26
xunit36-3  36  3  unitrc1  ra=5004.20  tb=0.05
xunit36-4  36  4  unitrc1  ra=1788.09  tb=0.06
xunit36-7  36  7  unitrc1  ra=8727.46  tb=0.04
xunit36-9  36  9  unitrc1  ra=2542.99  tb=0.08
xunit36-11  36  11  unitrc1  ra=7109.68  tb=0.04
xunit36-14  36  14  unitrc1  ra=4611.73  tb=0.46
xunit36-15  36  15  unitrc1  ra=1415.67  tb=0.13
xunit36-17  36  17  unitrc1  ra=9726.54  tb=0.35
xunit36-19  36  19  unitrc1  ra=5191.23  tb=0.32
xunit36-21  36  21  unitrc1  ra=9162.71  tb=0.48
xunit36-23  36  23  unitrc1  ra=1728.69  tb=0.06
xunit36-24  36  24  unitrc1  ra=2464.72  tb=0.13
xunit36-29  36  29  unitrc1  ra=3510.00  tb=0.36
xunit36-30  36  30  unitrc1  ra=1753.54  tb=0.35
xunit36-31  36  31  unitrc1  ra=638.32  tb=0.37
xunit36-32  36  32  unitrc1  ra=586.91  tb=0.23
xunit36-33  36  33  unitrc1  ra=7510.40  tb=0.38
xunit36-36  36  36  unitrc1  ra=2904.83  tb=0.09
xunit36-37  36  37  unitrc1  ra=4626.33  tb=0.05
xunit36-38  36  38  unitrc1  ra=2328.80  tb=0.07
xunit36-40  36  40  unitrc1  ra=6795.39  tb=0.16
xunit36-41  36  41  unitrc1  ra=4010.03  tb=0.20
xunit36-46  36  46  unitrc1  ra=4789.12  tb=0.29
xunit36-47  36  47  unitrc1  ra=294.97  tb=0.39

xunit37-5  37  5  unitrc1  ra=4908.86  tb=0.49
xunit37-6  37  6  unitrc1  ra=2168.71  tb=0.07
xunit37-10  37  10  unitrc1  ra=6644.03  tb=0.33
xunit37-11  37  11  unitrc1  ra=6273.21  tb=0.34
xunit37-12  37  12  unitrc1  ra=4786.90  tb=0.06
xunit37-14  37  14  unitrc1  ra=2106.77  tb=0.28
xunit37-16  37  16  unitrc1  ra=5048.29  tb=0.40
xunit37-18  37  18  unitrc1  ra=5106.93  tb=0.41
xunit37-19  37  19  unitrc1  ra=5849.22  tb=0.34
xunit37-20  37  20  unitrc1  ra=3288.12  tb=0.47
xunit37-21  37  21  unitrc1  ra=7553.70  tb=0.08
xunit37-23  37  23  unitrc1  ra=3370.78  tb=0.39
xunit37-24  37  24  unitrc1  ra=6657.02  tb=0.32
xunit37-25  37  25  unitrc1  ra=6595.72  tb=0.47
xunit37-26  37  26  unitrc1  ra=3876.19  tb=0.40
xunit37-28  37  28  unitrc1  ra=3373.40  tb=0.26
xunit37-29  37  29  unitrc1  ra=2804.13  tb=0.25
xunit37-30  37  30  unitrc1  ra=3720.04  tb=0.06
xunit37-32  37  32  unitrc1  ra=1795.13  tb=0.22
xunit37-33  37  33  unitrc1  ra=8987.97  tb=0.17
xunit37-34  37  34  unitrc1  ra=4052.12  tb=0.24
xunit37-36  37  36  unitrc1  ra=5297.11  tb=0.33
xunit37-37  37  37  unitrc1  ra=3979.69  tb=0.29
xunit37-38  37  38  unitrc1  ra=9290.06  tb=0.38
xunit37-39  37  39  unitrc1  ra=3672.06  tb=0.10
xunit37-41  37  41  unitrc1  ra=1489.25  tb=0.38
xunit37-42  37  42  unitrc1  ra=771.25  tb=0.44
xunit37-44  37  44  unitrc1  ra=3871.99  tb=0.37
xunit37-45  37  45  unitrc1  ra=7636.37  tb=0.25
xunit37-48  37  48  unitrc1  ra=3676.47  tb=0.21

xunit38-1  38  1  unitrc1  ra=4944.20  tb=0.07
xunit38-4  38  4  unitrc1  ra=6103.71  tb=0.26
xunit38-5  38  5  unitrc1  ra=2094.70  tb=0.21
xunit38-7  38  7  unitrc1  ra=9508.83  tb=0.04
xunit38-8  38  8  unitrc1  ra=2426.25  tb=0.41
xunit38-9  38  9  unitrc1  ra=7822.11  tb=0.19
xunit38-12  38  12  unitrc1  ra=4697.90  tb=0.06
xunit38-15  38  15  unitrc1  ra=7813.57  tb=0.26
xunit38-16  38  16  unitrc1  ra=4830.25  tb=0.03
xunit38-19  38  19  unitrc1  ra=4071.58  tb=0.29
xunit38-20  38  20  unitrc1  ra=6330.58  tb=0.00
xunit38-21  38  21  unitrc1  ra=9725.08  tb=0.33
xunit38-22  38  22  unitrc1  ra=3399.45  tb=0.33
xunit38-24  38  24  unitrc1  ra=7759.30  tb=0.22
xunit38-26  38  26  unitrc1  ra=1814.71  tb=0.17
xunit38-29  38  29  unitrc1  ra=3651.33  tb=0.15
xunit38-30  38  30  unitrc1  ra=5025.66  tb=0.40
xunit38-31  38  31  unitrc1  ra=400.91  tb=0.10
xunit38-32  38  32  unitrc1  ra=4462.85  tb=0.18
xunit38-35  38  35  unitrc1  ra=9596.48  tb=0.03
xunit38-37  38  37  unitrc1  ra=2990.54  tb=0.49
xunit38-38  38  38  unitrc1  ra=4534.97  tb=0.17
xunit38-39  38  39  unitrc1  ra=3783.34  tb=0.15
xunit38-40  38  40  unitrc1  ra=1809.84  tb=0.30
xunit38-42  38  42  unitrc1  ra=5011.57  tb=0.37
xunit38-47  38  47  unitrc1  ra=2329.03  tb=0.08
xunit38-48  38  48  unitrc1  ra=2818.92  tb=0.03
xunit38-49  38  49  unitrc1  ra=3415.96  tb=0.24
xunit38-50  38  50  unitrc1  ra=4525.51  tb=0.20

xunit39-1  39  1  unitrc1  ra=3171.64  tb=0.50
xunit39-2  39  2  unitrc1  ra=3507.35  tb=0.06
xunit39-3  39  3  unitrc1  ra=9688.07  tb=0.36
xunit39-5  39  5  unitrc1  ra=988.67  tb=0.41
xunit39-6  39  6  unitrc1  ra=6079.95  tb=0.28
xunit39-7  39  7  unitrc1  ra=2289.21  tb=0.30
xunit39-8  39  8  unitrc1  ra=6264.29  tb=0.26
xunit39-10  39  10  unitrc1  ra=7013.76  tb=0.17
xunit39-11  39  11  unitrc1  ra=1774.30  tb=0.03
xunit39-12  39  12  unitrc1  ra=5480.52  tb=0.17
xunit39-13  39  13  unitrc1  ra=9851.26  tb=0.26
xunit39-14  39  14  unitrc1  ra=4432.85  tb=0.48
xunit39-15  39  15  unitrc1  ra=862.75  tb=0.04
xunit39-16  39  16  unitrc1  ra=3993.19  tb=0.39
xunit39-18  39  18  unitrc1  ra=2323.62  tb=0.15
xunit39-22  39  22  unitrc1  ra=6518.69  tb=0.20
xunit39-23  39  23  unitrc1  ra=175.87  tb=0.02
xunit39-24  39  24  unitrc1  ra=5293.53  tb=0.17
xunit39-27  39  27  unitrc1  ra=6125.17  tb=0.40
xunit39-28  39  28  unitrc1  ra=7263.58  tb=0.08
xunit39-29  39  29  unitrc1  ra=3646.75  tb=0.10
xunit39-30  39  30  unitrc1  ra=3269.81  tb=0.19
xunit39-31  39  31  unitrc1  ra=7968.49  tb=0.08
xunit39-36  39  36  unitrc1  ra=1467.66  tb=0.40
xunit39-38  39  38  unitrc1  ra=413.97  tb=0.40
xunit39-39  39  39  unitrc1  ra=1116.26  tb=0.47
xunit39-40  39  40  unitrc1  ra=5842.30  tb=0.12
xunit39-43  39  43  unitrc1  ra=4955.50  tb=0.42
xunit39-45  39  45  unitrc1  ra=302.39  tb=0.31
xunit39-48  39  48  unitrc1  ra=225.77  tb=0.32
xunit39-49  39  49  unitrc1  ra=5577.44  tb=0.07

xunit40-2  40  2  unitrc1  ra=6111.43  tb=0.27
xunit40-4  40  4  unitrc1  ra=6670.77  tb=0.18
xunit40-5  40  5  unitrc1  ra=6603.74  tb=0.17
xunit40-8  40  8  unitrc1  ra=670.23  tb=0.49
xunit40-9  40  9  unitrc1  ra=311.55  tb=0.38
xunit40-10  40  10  unitrc1  ra=3985.98  tb=0.32
xunit40-11  40  11  unitrc1  ra=4588.44  tb=0.49
xunit40-12  40  12  unitrc1  ra=6622.97  tb=0.16
xunit40-14  40  14  unitrc1  ra=5047.96  tb=0.39
xunit40-17  40  17  unitrc1  ra=8054.89  tb=0.34
xunit40-18  40  18  unitrc1  ra=2443.74  tb=0.31
xunit40-19  40  19  unitrc1  ra=1224.55  tb=0.48
xunit40-21  40  21  unitrc1  ra=490.16  tb=0.04
xunit40-23  40  23  unitrc1  ra=3490.86  tb=0.42
xunit40-26  40  26  unitrc1  ra=6201.09  tb=0.39
xunit40-27  40  27  unitrc1  ra=2128.41  tb=0.43
xunit40-29  40  29  unitrc1  ra=3617.97  tb=0.28
xunit40-30  40  30  unitrc1  ra=3178.92  tb=0.40
xunit40-31  40  31  unitrc1  ra=4864.99  tb=0.30
xunit40-34  40  34  unitrc1  ra=961.14  tb=0.33
xunit40-35  40  35  unitrc1  ra=2587.78  tb=0.35
xunit40-36  40  36  unitrc1  ra=5449.47  tb=0.10
xunit40-39  40  39  unitrc1  ra=4626.94  tb=0.18
xunit40-40  40  40  unitrc1  ra=4839.98  tb=0.16
xunit40-41  40  41  unitrc1  ra=5927.96  tb=0.46
xunit40-42  40  42  unitrc1  ra=880.84  tb=0.29
xunit40-46  40  46  unitrc1  ra=7596.41  tb=0.25
xunit40-48  40  48  unitrc1  ra=1539.14  tb=0.13
xunit40-50  40  50  unitrc1  ra=7739.81  tb=0.30

xunit41-4  41  4  unitrc1  ra=830.18  tb=0.30
xunit41-5  41  5  unitrc1  ra=3362.97  tb=0.26
xunit41-6  41  6  unitrc1  ra=3064.45  tb=0.36
xunit41-7  41  7  unitrc1  ra=3969.33  tb=0.46
xunit41-11  41  11  unitrc1  ra=7169.95  tb=0.25
xunit41-15  41  15  unitrc1  ra=689.49  tb=0.20
xunit41-16  41  16  unitrc1  ra=2233.06  tb=0.15
xunit41-20  41  20  unitrc1  ra=1803.64  tb=0.21
xunit41-21  41  21  unitrc1  ra=2113.19  tb=0.09
xunit41-23  41  23  unitrc1  ra=8353.69  tb=0.11
xunit41-24  41  24  unitrc1  ra=3337.71  tb=0.26
xunit41-25  41  25  unitrc1  ra=2616.55  tb=0.28
xunit41-29  41  29  unitrc1  ra=7576.96  tb=0.30
xunit41-30  41  30  unitrc1  ra=3021.54  tb=0.09
xunit41-31  41  31  unitrc1  ra=1545.89  tb=0.50
xunit41-32  41  32  unitrc1  ra=5872.77  tb=0.38
xunit41-34  41  34  unitrc1  ra=2604.52  tb=0.45
xunit41-36  41  36  unitrc1  ra=7022.46  tb=0.39
xunit41-37  41  37  unitrc1  ra=2433.94  tb=0.36
xunit41-39  41  39  unitrc1  ra=3887.79  tb=0.47
xunit41-41  41  41  unitrc1  ra=6076.05  tb=0.32
xunit41-42  41  42  unitrc1  ra=1299.65  tb=0.12
xunit41-44  41  44  unitrc1  ra=5044.93  tb=0.25
xunit41-45  41  45  unitrc1  ra=6909.09  tb=0.32
xunit41-46  41  46  unitrc1  ra=2607.86  tb=0.38
xunit41-47  41  47  unitrc1  ra=3669.85  tb=0.41
xunit41-48  41  48  unitrc1  ra=4284.60  tb=0.31
xunit41-50  41  50  unitrc1  ra=5249.87  tb=0.15

xunit42-1  42  1  unitrc1  ra=3776.72  tb=0.34
xunit42-2  42  2  unitrc1  ra=3656.95  tb=0.22
xunit42-5  42  5  unitrc1  ra=3749.82  tb=0.03
xunit42-7  42  7  unitrc1  ra=3876.69  tb=0.42
xunit42-8  42  8  unitrc1  ra=9564.88  tb=0.09
xunit42-9  42  9  unitrc1  ra=8443.00  tb=0.29
xunit42-10  42  10  unitrc1  ra=7797.78  tb=0.31
xunit42-11  42  11  unitrc1  ra=8647.78  tb=0.11
xunit42-12  42  12  unitrc1  ra=1266.54  tb=0.04
xunit42-14  42  14  unitrc1  ra=2276.71  tb=0.19
xunit42-15  42  15  unitrc1  ra=5370.60  tb=0.37
xunit42-19  42  19  unitrc1  ra=805.75  tb=0.44
xunit42-21  42  21  unitrc1  ra=2008.88  tb=0.30
xunit42-22  42  22  unitrc1  ra=909.67  tb=0.42
xunit42-23  42  23  unitrc1  ra=8518.17  tb=0.20
xunit42-25  42  25  unitrc1  ra=4313.82  tb=0.28
xunit42-26  42  26  unitrc1  ra=5824.15  tb=0.09
xunit42-30  42  30  unitrc1  ra=9602.28  tb=0.48
xunit42-31  42  31  unitrc1  ra=3194.00  tb=0.48
xunit42-32  42  32  unitrc1  ra=4977.92  tb=0.31
xunit42-33  42  33  unitrc1  ra=6125.22  tb=0.16
xunit42-34  42  34  unitrc1  ra=508.34  tb=0.07
xunit42-35  42  35  unitrc1  ra=8710.07  tb=0.40
xunit42-36  42  36  unitrc1  ra=9220.71  tb=0.19
xunit42-37  42  37  unitrc1  ra=311.44  tb=0.41
xunit42-39  42  39  unitrc1  ra=4544.13  tb=0.33
xunit42-40  42  40  unitrc1  ra=7702.11  tb=0.21
xunit42-41  42  41  unitrc1  ra=5994.48  tb=0.29
xunit42-43  42  43  unitrc1  ra=5950.69  tb=0.38
xunit42-44  42  44  unitrc1  ra=7188.21  tb=0.16
xunit42-46  42  46  unitrc1  ra=9076.33  tb=0.40
xunit42-47  42  47  unitrc1  ra=3284.06  tb=0.37
xunit42-48  42  48  unitrc1  ra=9783.82  tb=0.27
xunit42-49  42  49  unitrc1  ra=6181.64  tb=0.04
xunit42-50  42  50  unitrc1  ra=2571.93  tb=0.43

xunit43-2  43  2  unitrc1  ra=4444.28  tb=0.09
xunit43-9  43  9  unitrc1  ra=3334.03  tb=0.26
xunit43-11  43  11  unitrc1  ra=3961.15  tb=0.03
xunit43-13  43  13  unitrc1  ra=4460.29  tb=0.03
xunit43-15  43  15  unitrc1  ra=8641.04  tb=0.20
xunit43-17  43  17  unitrc1  ra=708.23  tb=0.05
xunit43-20  43  20  unitrc1  ra=4471.81  tb=0.29
xunit43-21  43  21  unitrc1  ra=9571.79  tb=0.17
xunit43-22  43  22  unitrc1  ra=6885.47  tb=0.17
xunit43-23  43  23  unitrc1  ra=3315.73  tb=0.36
xunit43-26  43  26  unitrc1  ra=7420.40  tb=0.28
xunit43-28  43  28  unitrc1  ra=1128.46  tb=0.17
xunit43-29  43  29  unitrc1  ra=8296.00  tb=0.35
xunit43-32  43  32  unitrc1  ra=3096.69  tb=0.38
xunit43-33  43  33  unitrc1  ra=8405.11  tb=0.02
xunit43-36  43  36  unitrc1  ra=6382.87  tb=0.21
xunit43-39  43  39  unitrc1  ra=207.76  tb=0.13
xunit43-41  43  41  unitrc1  ra=6335.43  tb=0.20
xunit43-43  43  43  unitrc1  ra=9191.07  tb=0.14
xunit43-44  43  44  unitrc1  ra=7041.55  tb=0.23
xunit43-45  43  45  unitrc1  ra=2445.23  tb=0.43
xunit43-46  43  46  unitrc1  ra=4276.90  tb=0.04
xunit43-47  43  47  unitrc1  ra=3033.42  tb=0.35
xunit43-49  43  49  unitrc1  ra=1934.52  tb=0.12
xunit43-50  43  50  unitrc1  ra=4660.95  tb=0.32

xunit44-2  44  2  unitrc1  ra=3871.06  tb=0.37
xunit44-3  44  3  unitrc1  ra=4186.04  tb=0.32
xunit44-5  44  5  unitrc1  ra=7092.62  tb=0.09
xunit44-6  44  6  unitrc1  ra=2603.78  tb=0.45
xunit44-9  44  9  unitrc1  ra=322.02  tb=0.32
xunit44-10  44  10  unitrc1  ra=1099.43  tb=0.08
xunit44-11  44  11  unitrc1  ra=8035.48  tb=0.07
xunit44-12  44  12  unitrc1  ra=1984.81  tb=0.27
xunit44-13  44  13  unitrc1  ra=2090.84  tb=0.09
xunit44-14  44  14  unitrc1  ra=8354.06  tb=0.04
xunit44-15  44  15  unitrc1  ra=7463.52  tb=0.03
xunit44-16  44  16  unitrc1  ra=4366.09  tb=0.37
xunit44-17  44  17  unitrc1  ra=4050.80  tb=0.46
xunit44-19  44  19  unitrc1  ra=3288.44  tb=0.08
xunit44-21  44  21  unitrc1  ra=6990.23  tb=0.34
xunit44-23  44  23  unitrc1  ra=8479.57  tb=0.08
xunit44-25  44  25  unitrc1  ra=2001.25  tb=0.46
xunit44-28  44  28  unitrc1  ra=1463.02  tb=0.39
xunit44-32  44  32  unitrc1  ra=9499.99  tb=0.11
xunit44-35  44  35  unitrc1  ra=5036.39  tb=0.47
xunit44-38  44  38  unitrc1  ra=829.01  tb=0.45
xunit44-40  44  40  unitrc1  ra=8708.24  tb=0.32
xunit44-41  44  41  unitrc1  ra=3563.60  tb=0.28
xunit44-43  44  43  unitrc1  ra=1687.47  tb=0.45
xunit44-45  44  45  unitrc1  ra=9503.41  tb=0.23
xunit44-46  44  46  unitrc1  ra=9555.85  tb=0.20
xunit44-47  44  47  unitrc1  ra=3682.70  tb=0.47
xunit44-48  44  48  unitrc1  ra=8896.18  tb=0.16
xunit44-49  44  49  unitrc1  ra=7427.48  tb=0.18
xunit44-50  44  50  unitrc1  ra=3022.94  tb=0.21

xunit45-4  45  4  unitrc1  ra=3273.36  tb=0.11
xunit45-5  45  5  unitrc1  ra=4091.32  tb=0.02
xunit45-6  45  6  unitrc1  ra=5537.71  tb=0.23
xunit45-7  45  7  unitrc1  ra=6601.64  tb=0.09
xunit45-9  45  9  unitrc1  ra=6250.08  tb=0.05
xunit45-11  45  11  unitrc1  ra=3960.51  tb=0.18
xunit45-14  45  14  unitrc1  ra=3629.11  tb=0.36
xunit45-15  45  15  unitrc1  ra=1735.07  tb=0.43
xunit45-16  45  16  unitrc1  ra=2126.70  tb=0.03
xunit45-17  45  17  unitrc1  ra=153.82  tb=0.17
xunit45-18  45  18  unitrc1  ra=3444.45  tb=0.25
xunit45-19  45  19  unitrc1  ra=6670.95  tb=0.43
xunit45-21  45  21  unitrc1  ra=1379.22  tb=0.48
xunit45-22  45  22  unitrc1  ra=3396.50  tb=0.20
xunit45-23  45  23  unitrc1  ra=4203.21  tb=0.24
xunit45-25  45  25  unitrc1  ra=1274.13  tb=0.07
xunit45-26  45  26  unitrc1  ra=1683.24  tb=0.26
xunit45-27  45  27  unitrc1  ra=2149.03  tb=0.23
xunit45-28  45  28  unitrc1  ra=6583.10  tb=0.31
xunit45-29  45  29  unitrc1  ra=2019.92  tb=0.24
xunit45-30  45  30  unitrc1  ra=6705.67  tb=0.06
xunit45-31  45  31  unitrc1  ra=4458.09  tb=0.23
xunit45-32  45  32  unitrc1  ra=9451.50  tb=0.32
xunit45-37  45  37  unitrc1  ra=9037.38  tb=0.41
xunit45-38  45  38  unitrc1  ra=5962.07  tb=0.37
xunit45-39  45  39  unitrc1  ra=4846.48  tb=0.46
xunit45-40  45  40  unitrc1  ra=3970.87  tb=0.29
xunit45-43  45  43  unitrc1  ra=4703.14  tb=0.23
xunit45-44  45  44  unitrc1  ra=4150.41  tb=0.06
xunit45-45  45  45  unitrc1  ra=7664.23  tb=0.36
xunit45-46  45  46  unitrc1  ra=5272.48  tb=0.28
xunit45-47  45  47  unitrc1  ra=7853.71  tb=0.30
xunit45-49  45  49  unitrc1  ra=2328.40  tb=0.02

xunit46-2  46  2  unitrc1  ra=5621.07  tb=0.42
xunit46-6  46  6  unitrc1  ra=5264.16  tb=0.27
xunit46-7  46  7  unitrc1  ra=4744.72  tb=0.29
xunit46-13  46  13  unitrc1  ra=7908.59  tb=0.31
xunit46-14  46  14  unitrc1  ra=2640.12  tb=0.06
xunit46-17  46  17  unitrc1  ra=825.34  tb=0.44
xunit46-19  46  19  unitrc1  ra=3713.34  tb=0.48
xunit46-20  46  20  unitrc1  ra=9898.84  tb=0.20
xunit46-22  46  22  unitrc1  ra=7079.14  tb=0.12
xunit46-24  46  24  unitrc1  ra=4986.52  tb=0.50
xunit46-26  46  26  unitrc1  ra=2531.17  tb=0.11
xunit46-27  46  27  unitrc1  ra=7225.88  tb=0.30
xunit46-29  46  29  unitrc1  ra=2549.56  tb=0.47
xunit46-30  46  30  unitrc1  ra=2533.14  tb=0.48
xunit46-31  46  31  unitrc1  ra=3121.73  tb=0.49
xunit46-32  46  32  unitrc1  ra=9024.79  tb=0.37
xunit46-35  46  35  unitrc1  ra=1162.88  tb=0.35
xunit46-38  46  38  unitrc1  ra=3611.92  tb=0.14
xunit46-40  46  40  unitrc1  ra=1897.26  tb=0.16
xunit46-41  46  41  unitrc1  ra=4704.50  tb=0.46
xunit46-46  46  46  unitrc1  ra=6385.70  tb=0.46
xunit46-47  46  47  unitrc1  ra=2094.40  tb=0.46
xunit46-48  46  48  unitrc1  ra=7670.12  tb=0.14
xunit46-49  46  49  unitrc1  ra=1281.81  tb=0.30
xunit46-50  46  50  unitrc1  ra=1974.63  tb=0.22

xunit47-1  47  1  unitrc1  ra=6473.83  tb=0.03
xunit47-2  47  2  unitrc1  ra=7885.47  tb=0.42
xunit47-3  47  3  unitrc1  ra=5042.25  tb=0.13
xunit47-4  47  4  unitrc1  ra=748.84  tb=0.37
xunit47-5  47  5  unitrc1  ra=1620.50  tb=0.48
xunit47-6  47  6  unitrc1  ra=2591.55  tb=0.20
xunit47-7  47  7  unitrc1  ra=5860.45  tb=0.05
xunit47-9  47  9  unitrc1  ra=6318.96  tb=0.42
xunit47-11  47  11  unitrc1  ra=5721.29  tb=0.05
xunit47-13  47  13  unitrc1  ra=1430.49  tb=0.17
xunit47-14  47  14  unitrc1  ra=5347.31  tb=0.05
xunit47-19  47  19  unitrc1  ra=3635.63  tb=0.01
xunit47-20  47  20  unitrc1  ra=5736.80  tb=0.12
xunit47-21  47  21  unitrc1  ra=3101.73  tb=0.27
xunit47-22  47  22  unitrc1  ra=117.76  tb=0.02
xunit47-23  47  23  unitrc1  ra=5695.12  tb=0.39
xunit47-24  47  24  unitrc1  ra=6249.67  tb=0.31
xunit47-26  47  26  unitrc1  ra=3202.73  tb=0.19
xunit47-29  47  29  unitrc1  ra=5998.56  tb=0.36
xunit47-31  47  31  unitrc1  ra=5756.94  tb=0.27
xunit47-32  47  32  unitrc1  ra=810.45  tb=0.25
xunit47-33  47  33  unitrc1  ra=795.99  tb=0.03
xunit47-35  47  35  unitrc1  ra=3756.64  tb=0.19
xunit47-38  47  38  unitrc1  ra=5212.73  tb=0.16
xunit47-39  47  39  unitrc1  ra=2920.69  tb=0.09
xunit47-41  47  41  unitrc1  ra=3693.04  tb=0.37
xunit47-42  47  42  unitrc1  ra=6463.57  tb=0.39
xunit47-43  47  43  unitrc1  ra=3684.82  tb=0.14
xunit47-44  47  44  unitrc1  ra=4961.50  tb=0.17
xunit47-46  47  46  unitrc1  ra=6778.88  tb=0.23
xunit47-48  47  48  unitrc1  ra=728.45  tb=0.30
xunit47-50  47  50  unitrc1  ra=1507.28  tb=0.22

xunit48-3  48  3  unitrc1  ra=3880.97  tb=0.30
xunit48-5  48  5  unitrc1  ra=7963.61  tb=0.47
xunit48-7  48  7  unitrc1  ra=9278.78  tb=0.48
xunit48-9  48  9  unitrc1  ra=1339.95  tb=0.09
xunit48-11  48  11  unitrc1  ra=7537.20  tb=0.28
xunit48-12  48  12  unitrc1  ra=4272.46  tb=0.13
xunit48-13  48  13  unitrc1  ra=2606.18  tb=0.36
xunit48-14  48  14  unitrc1  ra=3893.51  tb=0.49
xunit48-17  48  17  unitrc1  ra=4805.32  tb=0.38
xunit48-18  48  18  unitrc1  ra=858.42  tb=0.35
xunit48-19  48  19  unitrc1  ra=1507.02  tb=0.25
xunit48-20  48  20  unitrc1  ra=7887.37  tb=0.36
xunit48-21  48  21  unitrc1  ra=3839.39  tb=0.46
xunit48-22  48  22  unitrc1  ra=8054.21  tb=0.49
xunit48-25  48  25  unitrc1  ra=9377.65  tb=0.40
xunit48-27  48  27  unitrc1  ra=5355.04  tb=0.45
xunit48-28  48  28  unitrc1  ra=139.09  tb=0.32
xunit48-30  48  30  unitrc1  ra=5693.99  tb=0.06
xunit48-31  48  31  unitrc1  ra=3220.52  tb=0.22
xunit48-33  48  33  unitrc1  ra=1903.20  tb=0.07
xunit48-36  48  36  unitrc1  ra=6404.48  tb=0.22
xunit48-37  48  37  unitrc1  ra=611.76  tb=0.36
xunit48-38  48  38  unitrc1  ra=6832.67  tb=0.01
xunit48-40  48  40  unitrc1  ra=3844.30  tb=0.35
xunit48-41  48  41  unitrc1  ra=3439.27  tb=0.24
xunit48-42  48  42  unitrc1  ra=8308.26  tb=0.18
xunit48-45  48  45  unitrc1  ra=3263.39  tb=0.25
xunit48-49  48  49  unitrc1  ra=4209.20  tb=0.28

xunit49-2  49  2  unitrc1  ra=7528.02  tb=0.26
xunit49-3  49  3  unitrc1  ra=6613.43  tb=0.10
xunit49-6  49  6  unitrc1  ra=3947.53  tb=0.09
xunit49-7  49  7  unitrc1  ra=357.40  tb=0.45
xunit49-8  49  8  unitrc1  ra=5312.33  tb=0.07
xunit49-9  49  9  unitrc1  ra=5423.98  tb=0.31
xunit49-10  49  10  unitrc1  ra=4156.33  tb=0.01
xunit49-11  49  11  unitrc1  ra=2394.74  tb=0.42
xunit49-12  49  12  unitrc1  ra=350.56  tb=0.43
xunit49-15  49  15  unitrc1  ra=6067.51  tb=0.45
xunit49-16  49  16  unitrc1  ra=7182.16  tb=0.21
xunit49-17  49  17  unitrc1  ra=2533.83  tb=0.34
xunit49-18  49  18  unitrc1  ra=8713.16  tb=0.26
xunit49-22  49  22  unitrc1  ra=9193.31  tb=0.01
xunit49-23  49  23  unitrc1  ra=1881.19  tb=0.37
xunit49-24  49  24  unitrc1  ra=7264.27  tb=0.25
xunit49-25  49  25  unitrc1  ra=6016.29  tb=0.20
xunit49-27  49  27  unitrc1  ra=5331.73  tb=0.09
xunit49-29  49  29  unitrc1  ra=1804.45  tb=0.05
xunit49-30  49  30  unitrc1  ra=2706.58  tb=0.24
xunit49-31  49  31  unitrc1  ra=6622.68  tb=0.41
xunit49-33  49  33  unitrc1  ra=3220.55  tb=0.15
xunit49-34  49  34  unitrc1  ra=3370.38  tb=0.01
xunit49-37  49  37  unitrc1  ra=4253.61  tb=0.15
xunit49-39  49  39  unitrc1  ra=6242.20  tb=0.39
xunit49-41  49  41  unitrc1  ra=2456.77  tb=0.11
xunit49-42  49  42  unitrc1  ra=368.02  tb=0.38
xunit49-43  49  43  unitrc1  ra=8277.12  tb=0.22
xunit49-45  49  45  unitrc1  ra=2212.67  tb=0.20
xunit49-46  49  46  unitrc1  ra=6271.46  tb=0.29
xunit49-47  49  47  unitrc1  ra=5905.36  tb=0.45
xunit49-48  49  48  unitrc1  ra=7962.45  tb=0.02
xunit49-49  49  49  unitrc1  ra=3407.95  tb=0.11
xunit49-50  49  50  unitrc1  ra=8549.79  tb=0.20

xunit50-4  50  4  unitrc1  ra=2511.94  tb=0.28
xunit50-5  50  5  unitrc1  ra=842.40  tb=0.21
xunit50-6  50  6  unitrc1  ra=2103.71  tb=0.34
xunit50-7  50  7  unitrc1  ra=8117.20  tb=0.42
xunit50-8  50  8  unitrc1  ra=2170.83  tb=0.33
xunit50-9  50  9  unitrc1  ra=3573.49  tb=0.50
xunit50-11  50  11  unitrc1  ra=6361.91  tb=0.13
xunit50-13  50  13  unitrc1  ra=1825.81  tb=0.09
xunit50-15  50  15  unitrc1  ra=5221.20  tb=0.30
xunit50-16  50  16  unitrc1  ra=4041.83  tb=0.01
xunit50-17  50  17  unitrc1  ra=2614.81  tb=0.42
xunit50-18  50  18  unitrc1  ra=9360.96  tb=0.34
xunit50-19  50  19  unitrc1  ra=9171.42  tb=0.22
xunit50-20  50  20  unitrc1  ra=219.79  tb=0.44
xunit50-21  50  21  unitrc1  ra=7691.26  tb=0.32
xunit50-24  50  24  unitrc1  ra=662.63  tb=0.03
xunit50-25  50  25  unitrc1  ra=7125.67  tb=0.43
xunit50-27  50  27  unitrc1  ra=6477.32  tb=0.07
xunit50-28  50  28  unitrc1  ra=6882.75  tb=0.12
xunit50-29  50  29  unitrc1  ra=4842.28  tb=0.19
xunit50-30  50  30  unitrc1  ra=6505.75  tb=0.31
xunit50-32  50  32  unitrc1  ra=7448.62  tb=0.00
xunit50-33  50  33  unitrc1  ra=2344.64  tb=0.11
xunit50-34  50  34  unitrc1  ra=3949.10  tb=0.43
xunit50-35  50  35  unitrc1  ra=822.82  tb=0.32
xunit50-37  50  37  unitrc1  ra=5379.70  tb=0.44
xunit50-39  50  39  unitrc1  ra=5920.08  tb=0.08
xunit50-44  50  44  unitrc1  ra=5508.02  tb=0.46
xunit50-46  50  46  unitrc1  ra=7808.43  tb=0.30
xunit50-47  50  47  unitrc1  ra=1873.06  tb=0.46
xunit50-48  50  48  unitrc1  ra=3531.41  tb=0.24
xunit50-49  50  49  unitrc1  ra=3487.14  tb=0.08

.save   time
.save   v.xunit1-1.vtemp2#branch
.save   v.xunit1-2.vtemp2#branch
.save   v.xunit1-3.vtemp2#branch
.save   v.xunit1-4.vtemp2#branch
.save   v.xunit1-5.vtemp2#branch
.save   v.xunit1-6.vtemp2#branch
.save   v.xunit1-7.vtemp2#branch
.save   v.xunit1-8.vtemp2#branch
.save   v.xunit1-9.vtemp2#branch
.save   v.xunit1-10.vtemp2#branch
.save   v.xunit1-11.vtemp2#branch
.save   v.xunit1-12.vtemp2#branch
.save   v.xunit1-13.vtemp2#branch
.save   v.xunit1-14.vtemp2#branch
.save   v.xunit1-15.vtemp2#branch
.save   v.xunit1-16.vtemp2#branch
.save   v.xunit1-17.vtemp2#branch
.save   v.xunit1-18.vtemp2#branch
.save   v.xunit1-19.vtemp2#branch
.save   v.xunit1-20.vtemp2#branch
.save   v.xunit1-21.vtemp2#branch
.save   v.xunit1-22.vtemp2#branch
.save   v.xunit1-23.vtemp2#branch
.save   v.xunit1-24.vtemp2#branch
.save   v.xunit1-25.vtemp2#branch
.save   v.xunit1-26.vtemp2#branch
.save   v.xunit1-27.vtemp2#branch
.save   v.xunit1-28.vtemp2#branch
.save   v.xunit1-29.vtemp2#branch
.save   v.xunit1-30.vtemp2#branch
.save   v.xunit1-31.vtemp2#branch
.save   v.xunit1-32.vtemp2#branch
.save   v.xunit1-33.vtemp2#branch
.save   v.xunit1-34.vtemp2#branch
.save   v.xunit1-35.vtemp2#branch
.save   v.xunit1-36.vtemp2#branch
.save   v.xunit1-37.vtemp2#branch
.save   v.xunit1-38.vtemp2#branch
.save   v.xunit1-39.vtemp2#branch
.save   v.xunit1-40.vtemp2#branch
.save   v.xunit1-41.vtemp2#branch
.save   v.xunit1-42.vtemp2#branch
.save   v.xunit1-43.vtemp2#branch
.save   v.xunit1-44.vtemp2#branch
.save   v.xunit1-45.vtemp2#branch
.save   v.xunit1-46.vtemp2#branch
.save   v.xunit1-47.vtemp2#branch
.save   v.xunit1-48.vtemp2#branch
.save   v.xunit1-49.vtemp2#branch
.save   v.xunit1-50.vtemp2#branch

.save   v.xunit2-1.vtemp2#branch
.save   v.xunit2-2.vtemp2#branch
.save   v.xunit2-3.vtemp2#branch
.save   v.xunit2-4.vtemp2#branch
.save   v.xunit2-5.vtemp2#branch
.save   v.xunit2-6.vtemp2#branch
.save   v.xunit2-7.vtemp2#branch
.save   v.xunit2-8.vtemp2#branch
.save   v.xunit2-9.vtemp2#branch
.save   v.xunit2-10.vtemp2#branch
.save   v.xunit2-11.vtemp2#branch
.save   v.xunit2-12.vtemp2#branch
.save   v.xunit2-13.vtemp2#branch
.save   v.xunit2-14.vtemp2#branch
.save   v.xunit2-15.vtemp2#branch
.save   v.xunit2-16.vtemp2#branch
.save   v.xunit2-17.vtemp2#branch
.save   v.xunit2-18.vtemp2#branch
.save   v.xunit2-19.vtemp2#branch
.save   v.xunit2-20.vtemp2#branch
.save   v.xunit2-21.vtemp2#branch
.save   v.xunit2-22.vtemp2#branch
.save   v.xunit2-23.vtemp2#branch
.save   v.xunit2-24.vtemp2#branch
.save   v.xunit2-25.vtemp2#branch
.save   v.xunit2-26.vtemp2#branch
.save   v.xunit2-27.vtemp2#branch
.save   v.xunit2-28.vtemp2#branch
.save   v.xunit2-29.vtemp2#branch
.save   v.xunit2-30.vtemp2#branch
.save   v.xunit2-31.vtemp2#branch
.save   v.xunit2-32.vtemp2#branch
.save   v.xunit2-33.vtemp2#branch
.save   v.xunit2-34.vtemp2#branch
.save   v.xunit2-35.vtemp2#branch
.save   v.xunit2-36.vtemp2#branch
.save   v.xunit2-37.vtemp2#branch
.save   v.xunit2-38.vtemp2#branch
.save   v.xunit2-39.vtemp2#branch
.save   v.xunit2-40.vtemp2#branch
.save   v.xunit2-41.vtemp2#branch
.save   v.xunit2-42.vtemp2#branch
.save   v.xunit2-43.vtemp2#branch
.save   v.xunit2-44.vtemp2#branch
.save   v.xunit2-45.vtemp2#branch
.save   v.xunit2-46.vtemp2#branch
.save   v.xunit2-47.vtemp2#branch
.save   v.xunit2-48.vtemp2#branch
.save   v.xunit2-49.vtemp2#branch
.save   v.xunit2-50.vtemp2#branch

.save   v.xunit3-1.vtemp2#branch
.save   v.xunit3-2.vtemp2#branch
.save   v.xunit3-3.vtemp2#branch
.save   v.xunit3-4.vtemp2#branch
.save   v.xunit3-5.vtemp2#branch
.save   v.xunit3-6.vtemp2#branch
.save   v.xunit3-7.vtemp2#branch
.save   v.xunit3-8.vtemp2#branch
.save   v.xunit3-9.vtemp2#branch
.save   v.xunit3-10.vtemp2#branch
.save   v.xunit3-11.vtemp2#branch
.save   v.xunit3-12.vtemp2#branch
.save   v.xunit3-13.vtemp2#branch
.save   v.xunit3-14.vtemp2#branch
.save   v.xunit3-15.vtemp2#branch
.save   v.xunit3-16.vtemp2#branch
.save   v.xunit3-17.vtemp2#branch
.save   v.xunit3-18.vtemp2#branch
.save   v.xunit3-19.vtemp2#branch
.save   v.xunit3-20.vtemp2#branch
.save   v.xunit3-21.vtemp2#branch
.save   v.xunit3-22.vtemp2#branch
.save   v.xunit3-23.vtemp2#branch
.save   v.xunit3-24.vtemp2#branch
.save   v.xunit3-25.vtemp2#branch
.save   v.xunit3-26.vtemp2#branch
.save   v.xunit3-27.vtemp2#branch
.save   v.xunit3-28.vtemp2#branch
.save   v.xunit3-29.vtemp2#branch
.save   v.xunit3-30.vtemp2#branch
.save   v.xunit3-31.vtemp2#branch
.save   v.xunit3-32.vtemp2#branch
.save   v.xunit3-33.vtemp2#branch
.save   v.xunit3-34.vtemp2#branch
.save   v.xunit3-35.vtemp2#branch
.save   v.xunit3-36.vtemp2#branch
.save   v.xunit3-37.vtemp2#branch
.save   v.xunit3-38.vtemp2#branch
.save   v.xunit3-39.vtemp2#branch
.save   v.xunit3-40.vtemp2#branch
.save   v.xunit3-41.vtemp2#branch
.save   v.xunit3-42.vtemp2#branch
.save   v.xunit3-43.vtemp2#branch
.save   v.xunit3-44.vtemp2#branch
.save   v.xunit3-45.vtemp2#branch
.save   v.xunit3-46.vtemp2#branch
.save   v.xunit3-47.vtemp2#branch
.save   v.xunit3-48.vtemp2#branch
.save   v.xunit3-49.vtemp2#branch
.save   v.xunit3-50.vtemp2#branch

.save   v.xunit4-1.vtemp2#branch
.save   v.xunit4-2.vtemp2#branch
.save   v.xunit4-3.vtemp2#branch
.save   v.xunit4-4.vtemp2#branch
.save   v.xunit4-5.vtemp2#branch
.save   v.xunit4-6.vtemp2#branch
.save   v.xunit4-7.vtemp2#branch
.save   v.xunit4-8.vtemp2#branch
.save   v.xunit4-9.vtemp2#branch
.save   v.xunit4-10.vtemp2#branch
.save   v.xunit4-11.vtemp2#branch
.save   v.xunit4-12.vtemp2#branch
.save   v.xunit4-13.vtemp2#branch
.save   v.xunit4-14.vtemp2#branch
.save   v.xunit4-15.vtemp2#branch
.save   v.xunit4-16.vtemp2#branch
.save   v.xunit4-17.vtemp2#branch
.save   v.xunit4-18.vtemp2#branch
.save   v.xunit4-19.vtemp2#branch
.save   v.xunit4-20.vtemp2#branch
.save   v.xunit4-21.vtemp2#branch
.save   v.xunit4-22.vtemp2#branch
.save   v.xunit4-23.vtemp2#branch
.save   v.xunit4-24.vtemp2#branch
.save   v.xunit4-25.vtemp2#branch
.save   v.xunit4-26.vtemp2#branch
.save   v.xunit4-27.vtemp2#branch
.save   v.xunit4-28.vtemp2#branch
.save   v.xunit4-29.vtemp2#branch
.save   v.xunit4-30.vtemp2#branch
.save   v.xunit4-31.vtemp2#branch
.save   v.xunit4-32.vtemp2#branch
.save   v.xunit4-33.vtemp2#branch
.save   v.xunit4-34.vtemp2#branch
.save   v.xunit4-35.vtemp2#branch
.save   v.xunit4-36.vtemp2#branch
.save   v.xunit4-37.vtemp2#branch
.save   v.xunit4-38.vtemp2#branch
.save   v.xunit4-39.vtemp2#branch
.save   v.xunit4-40.vtemp2#branch
.save   v.xunit4-41.vtemp2#branch
.save   v.xunit4-42.vtemp2#branch
.save   v.xunit4-43.vtemp2#branch
.save   v.xunit4-44.vtemp2#branch
.save   v.xunit4-45.vtemp2#branch
.save   v.xunit4-46.vtemp2#branch
.save   v.xunit4-47.vtemp2#branch
.save   v.xunit4-48.vtemp2#branch
.save   v.xunit4-49.vtemp2#branch
.save   v.xunit4-50.vtemp2#branch

.save   v.xunit5-1.vtemp2#branch
.save   v.xunit5-2.vtemp2#branch
.save   v.xunit5-3.vtemp2#branch
.save   v.xunit5-4.vtemp2#branch
.save   v.xunit5-5.vtemp2#branch
.save   v.xunit5-6.vtemp2#branch
.save   v.xunit5-7.vtemp2#branch
.save   v.xunit5-8.vtemp2#branch
.save   v.xunit5-9.vtemp2#branch
.save   v.xunit5-10.vtemp2#branch
.save   v.xunit5-11.vtemp2#branch
.save   v.xunit5-12.vtemp2#branch
.save   v.xunit5-13.vtemp2#branch
.save   v.xunit5-14.vtemp2#branch
.save   v.xunit5-15.vtemp2#branch
.save   v.xunit5-16.vtemp2#branch
.save   v.xunit5-17.vtemp2#branch
.save   v.xunit5-18.vtemp2#branch
.save   v.xunit5-19.vtemp2#branch
.save   v.xunit5-20.vtemp2#branch
.save   v.xunit5-21.vtemp2#branch
.save   v.xunit5-22.vtemp2#branch
.save   v.xunit5-23.vtemp2#branch
.save   v.xunit5-24.vtemp2#branch
.save   v.xunit5-25.vtemp2#branch
.save   v.xunit5-26.vtemp2#branch
.save   v.xunit5-27.vtemp2#branch
.save   v.xunit5-28.vtemp2#branch
.save   v.xunit5-29.vtemp2#branch
.save   v.xunit5-30.vtemp2#branch
.save   v.xunit5-31.vtemp2#branch
.save   v.xunit5-32.vtemp2#branch
.save   v.xunit5-33.vtemp2#branch
.save   v.xunit5-34.vtemp2#branch
.save   v.xunit5-35.vtemp2#branch
.save   v.xunit5-36.vtemp2#branch
.save   v.xunit5-37.vtemp2#branch
.save   v.xunit5-38.vtemp2#branch
.save   v.xunit5-39.vtemp2#branch
.save   v.xunit5-40.vtemp2#branch
.save   v.xunit5-41.vtemp2#branch
.save   v.xunit5-42.vtemp2#branch
.save   v.xunit5-43.vtemp2#branch
.save   v.xunit5-44.vtemp2#branch
.save   v.xunit5-45.vtemp2#branch
.save   v.xunit5-46.vtemp2#branch
.save   v.xunit5-47.vtemp2#branch
.save   v.xunit5-48.vtemp2#branch
.save   v.xunit5-49.vtemp2#branch
.save   v.xunit5-50.vtemp2#branch

.save   v.xunit6-1.vtemp2#branch
.save   v.xunit6-2.vtemp2#branch
.save   v.xunit6-3.vtemp2#branch
.save   v.xunit6-4.vtemp2#branch
.save   v.xunit6-5.vtemp2#branch
.save   v.xunit6-6.vtemp2#branch
.save   v.xunit6-7.vtemp2#branch
.save   v.xunit6-8.vtemp2#branch
.save   v.xunit6-9.vtemp2#branch
.save   v.xunit6-10.vtemp2#branch
.save   v.xunit6-11.vtemp2#branch
.save   v.xunit6-12.vtemp2#branch
.save   v.xunit6-13.vtemp2#branch
.save   v.xunit6-14.vtemp2#branch
.save   v.xunit6-15.vtemp2#branch
.save   v.xunit6-16.vtemp2#branch
.save   v.xunit6-17.vtemp2#branch
.save   v.xunit6-18.vtemp2#branch
.save   v.xunit6-19.vtemp2#branch
.save   v.xunit6-20.vtemp2#branch
.save   v.xunit6-21.vtemp2#branch
.save   v.xunit6-22.vtemp2#branch
.save   v.xunit6-23.vtemp2#branch
.save   v.xunit6-24.vtemp2#branch
.save   v.xunit6-25.vtemp2#branch
.save   v.xunit6-26.vtemp2#branch
.save   v.xunit6-27.vtemp2#branch
.save   v.xunit6-28.vtemp2#branch
.save   v.xunit6-29.vtemp2#branch
.save   v.xunit6-30.vtemp2#branch
.save   v.xunit6-31.vtemp2#branch
.save   v.xunit6-32.vtemp2#branch
.save   v.xunit6-33.vtemp2#branch
.save   v.xunit6-34.vtemp2#branch
.save   v.xunit6-35.vtemp2#branch
.save   v.xunit6-36.vtemp2#branch
.save   v.xunit6-37.vtemp2#branch
.save   v.xunit6-38.vtemp2#branch
.save   v.xunit6-39.vtemp2#branch
.save   v.xunit6-40.vtemp2#branch
.save   v.xunit6-41.vtemp2#branch
.save   v.xunit6-42.vtemp2#branch
.save   v.xunit6-43.vtemp2#branch
.save   v.xunit6-44.vtemp2#branch
.save   v.xunit6-45.vtemp2#branch
.save   v.xunit6-46.vtemp2#branch
.save   v.xunit6-47.vtemp2#branch
.save   v.xunit6-48.vtemp2#branch
.save   v.xunit6-49.vtemp2#branch
.save   v.xunit6-50.vtemp2#branch

.save   v.xunit7-1.vtemp2#branch
.save   v.xunit7-2.vtemp2#branch
.save   v.xunit7-3.vtemp2#branch
.save   v.xunit7-4.vtemp2#branch
.save   v.xunit7-5.vtemp2#branch
.save   v.xunit7-6.vtemp2#branch
.save   v.xunit7-7.vtemp2#branch
.save   v.xunit7-8.vtemp2#branch
.save   v.xunit7-9.vtemp2#branch
.save   v.xunit7-10.vtemp2#branch
.save   v.xunit7-11.vtemp2#branch
.save   v.xunit7-12.vtemp2#branch
.save   v.xunit7-13.vtemp2#branch
.save   v.xunit7-14.vtemp2#branch
.save   v.xunit7-15.vtemp2#branch
.save   v.xunit7-16.vtemp2#branch
.save   v.xunit7-17.vtemp2#branch
.save   v.xunit7-18.vtemp2#branch
.save   v.xunit7-19.vtemp2#branch
.save   v.xunit7-20.vtemp2#branch
.save   v.xunit7-21.vtemp2#branch
.save   v.xunit7-22.vtemp2#branch
.save   v.xunit7-23.vtemp2#branch
.save   v.xunit7-24.vtemp2#branch
.save   v.xunit7-25.vtemp2#branch
.save   v.xunit7-26.vtemp2#branch
.save   v.xunit7-27.vtemp2#branch
.save   v.xunit7-28.vtemp2#branch
.save   v.xunit7-29.vtemp2#branch
.save   v.xunit7-30.vtemp2#branch
.save   v.xunit7-31.vtemp2#branch
.save   v.xunit7-32.vtemp2#branch
.save   v.xunit7-33.vtemp2#branch
.save   v.xunit7-34.vtemp2#branch
.save   v.xunit7-35.vtemp2#branch
.save   v.xunit7-36.vtemp2#branch
.save   v.xunit7-37.vtemp2#branch
.save   v.xunit7-38.vtemp2#branch
.save   v.xunit7-39.vtemp2#branch
.save   v.xunit7-40.vtemp2#branch
.save   v.xunit7-41.vtemp2#branch
.save   v.xunit7-42.vtemp2#branch
.save   v.xunit7-43.vtemp2#branch
.save   v.xunit7-44.vtemp2#branch
.save   v.xunit7-45.vtemp2#branch
.save   v.xunit7-46.vtemp2#branch
.save   v.xunit7-47.vtemp2#branch
.save   v.xunit7-48.vtemp2#branch
.save   v.xunit7-49.vtemp2#branch
.save   v.xunit7-50.vtemp2#branch

.save   v.xunit8-1.vtemp2#branch
.save   v.xunit8-2.vtemp2#branch
.save   v.xunit8-3.vtemp2#branch
.save   v.xunit8-4.vtemp2#branch
.save   v.xunit8-5.vtemp2#branch
.save   v.xunit8-6.vtemp2#branch
.save   v.xunit8-7.vtemp2#branch
.save   v.xunit8-8.vtemp2#branch
.save   v.xunit8-9.vtemp2#branch
.save   v.xunit8-10.vtemp2#branch
.save   v.xunit8-11.vtemp2#branch
.save   v.xunit8-12.vtemp2#branch
.save   v.xunit8-13.vtemp2#branch
.save   v.xunit8-14.vtemp2#branch
.save   v.xunit8-15.vtemp2#branch
.save   v.xunit8-16.vtemp2#branch
.save   v.xunit8-17.vtemp2#branch
.save   v.xunit8-18.vtemp2#branch
.save   v.xunit8-19.vtemp2#branch
.save   v.xunit8-20.vtemp2#branch
.save   v.xunit8-21.vtemp2#branch
.save   v.xunit8-22.vtemp2#branch
.save   v.xunit8-23.vtemp2#branch
.save   v.xunit8-24.vtemp2#branch
.save   v.xunit8-25.vtemp2#branch
.save   v.xunit8-26.vtemp2#branch
.save   v.xunit8-27.vtemp2#branch
.save   v.xunit8-28.vtemp2#branch
.save   v.xunit8-29.vtemp2#branch
.save   v.xunit8-30.vtemp2#branch
.save   v.xunit8-31.vtemp2#branch
.save   v.xunit8-32.vtemp2#branch
.save   v.xunit8-33.vtemp2#branch
.save   v.xunit8-34.vtemp2#branch
.save   v.xunit8-35.vtemp2#branch
.save   v.xunit8-36.vtemp2#branch
.save   v.xunit8-37.vtemp2#branch
.save   v.xunit8-38.vtemp2#branch
.save   v.xunit8-39.vtemp2#branch
.save   v.xunit8-40.vtemp2#branch
.save   v.xunit8-41.vtemp2#branch
.save   v.xunit8-42.vtemp2#branch
.save   v.xunit8-43.vtemp2#branch
.save   v.xunit8-44.vtemp2#branch
.save   v.xunit8-45.vtemp2#branch
.save   v.xunit8-46.vtemp2#branch
.save   v.xunit8-47.vtemp2#branch
.save   v.xunit8-48.vtemp2#branch
.save   v.xunit8-49.vtemp2#branch
.save   v.xunit8-50.vtemp2#branch

.save   v.xunit9-1.vtemp2#branch
.save   v.xunit9-2.vtemp2#branch
.save   v.xunit9-3.vtemp2#branch
.save   v.xunit9-4.vtemp2#branch
.save   v.xunit9-5.vtemp2#branch
.save   v.xunit9-6.vtemp2#branch
.save   v.xunit9-7.vtemp2#branch
.save   v.xunit9-8.vtemp2#branch
.save   v.xunit9-9.vtemp2#branch
.save   v.xunit9-10.vtemp2#branch
.save   v.xunit9-11.vtemp2#branch
.save   v.xunit9-12.vtemp2#branch
.save   v.xunit9-13.vtemp2#branch
.save   v.xunit9-14.vtemp2#branch
.save   v.xunit9-15.vtemp2#branch
.save   v.xunit9-16.vtemp2#branch
.save   v.xunit9-17.vtemp2#branch
.save   v.xunit9-18.vtemp2#branch
.save   v.xunit9-19.vtemp2#branch
.save   v.xunit9-20.vtemp2#branch
.save   v.xunit9-21.vtemp2#branch
.save   v.xunit9-22.vtemp2#branch
.save   v.xunit9-23.vtemp2#branch
.save   v.xunit9-24.vtemp2#branch
.save   v.xunit9-25.vtemp2#branch
.save   v.xunit9-26.vtemp2#branch
.save   v.xunit9-27.vtemp2#branch
.save   v.xunit9-28.vtemp2#branch
.save   v.xunit9-29.vtemp2#branch
.save   v.xunit9-30.vtemp2#branch
.save   v.xunit9-31.vtemp2#branch
.save   v.xunit9-32.vtemp2#branch
.save   v.xunit9-33.vtemp2#branch
.save   v.xunit9-34.vtemp2#branch
.save   v.xunit9-35.vtemp2#branch
.save   v.xunit9-36.vtemp2#branch
.save   v.xunit9-37.vtemp2#branch
.save   v.xunit9-38.vtemp2#branch
.save   v.xunit9-39.vtemp2#branch
.save   v.xunit9-40.vtemp2#branch
.save   v.xunit9-41.vtemp2#branch
.save   v.xunit9-42.vtemp2#branch
.save   v.xunit9-43.vtemp2#branch
.save   v.xunit9-44.vtemp2#branch
.save   v.xunit9-45.vtemp2#branch
.save   v.xunit9-46.vtemp2#branch
.save   v.xunit9-47.vtemp2#branch
.save   v.xunit9-48.vtemp2#branch
.save   v.xunit9-49.vtemp2#branch
.save   v.xunit9-50.vtemp2#branch

.save   v.xunit10-1.vtemp2#branch
.save   v.xunit10-2.vtemp2#branch
.save   v.xunit10-3.vtemp2#branch
.save   v.xunit10-4.vtemp2#branch
.save   v.xunit10-5.vtemp2#branch
.save   v.xunit10-6.vtemp2#branch
.save   v.xunit10-7.vtemp2#branch
.save   v.xunit10-8.vtemp2#branch
.save   v.xunit10-9.vtemp2#branch
.save   v.xunit10-10.vtemp2#branch
.save   v.xunit10-11.vtemp2#branch
.save   v.xunit10-12.vtemp2#branch
.save   v.xunit10-13.vtemp2#branch
.save   v.xunit10-14.vtemp2#branch
.save   v.xunit10-15.vtemp2#branch
.save   v.xunit10-16.vtemp2#branch
.save   v.xunit10-17.vtemp2#branch
.save   v.xunit10-18.vtemp2#branch
.save   v.xunit10-19.vtemp2#branch
.save   v.xunit10-20.vtemp2#branch
.save   v.xunit10-21.vtemp2#branch
.save   v.xunit10-22.vtemp2#branch
.save   v.xunit10-23.vtemp2#branch
.save   v.xunit10-24.vtemp2#branch
.save   v.xunit10-25.vtemp2#branch
.save   v.xunit10-26.vtemp2#branch
.save   v.xunit10-27.vtemp2#branch
.save   v.xunit10-28.vtemp2#branch
.save   v.xunit10-29.vtemp2#branch
.save   v.xunit10-30.vtemp2#branch
.save   v.xunit10-31.vtemp2#branch
.save   v.xunit10-32.vtemp2#branch
.save   v.xunit10-33.vtemp2#branch
.save   v.xunit10-34.vtemp2#branch
.save   v.xunit10-35.vtemp2#branch
.save   v.xunit10-36.vtemp2#branch
.save   v.xunit10-37.vtemp2#branch
.save   v.xunit10-38.vtemp2#branch
.save   v.xunit10-39.vtemp2#branch
.save   v.xunit10-40.vtemp2#branch
.save   v.xunit10-41.vtemp2#branch
.save   v.xunit10-42.vtemp2#branch
.save   v.xunit10-43.vtemp2#branch
.save   v.xunit10-44.vtemp2#branch
.save   v.xunit10-45.vtemp2#branch
.save   v.xunit10-46.vtemp2#branch
.save   v.xunit10-47.vtemp2#branch
.save   v.xunit10-48.vtemp2#branch
.save   v.xunit10-49.vtemp2#branch
.save   v.xunit10-50.vtemp2#branch

.save   v.xunit11-1.vtemp2#branch
.save   v.xunit11-2.vtemp2#branch
.save   v.xunit11-3.vtemp2#branch
.save   v.xunit11-4.vtemp2#branch
.save   v.xunit11-5.vtemp2#branch
.save   v.xunit11-6.vtemp2#branch
.save   v.xunit11-7.vtemp2#branch
.save   v.xunit11-8.vtemp2#branch
.save   v.xunit11-9.vtemp2#branch
.save   v.xunit11-10.vtemp2#branch
.save   v.xunit11-11.vtemp2#branch
.save   v.xunit11-12.vtemp2#branch
.save   v.xunit11-13.vtemp2#branch
.save   v.xunit11-14.vtemp2#branch
.save   v.xunit11-15.vtemp2#branch
.save   v.xunit11-16.vtemp2#branch
.save   v.xunit11-17.vtemp2#branch
.save   v.xunit11-18.vtemp2#branch
.save   v.xunit11-19.vtemp2#branch
.save   v.xunit11-20.vtemp2#branch
.save   v.xunit11-21.vtemp2#branch
.save   v.xunit11-22.vtemp2#branch
.save   v.xunit11-23.vtemp2#branch
.save   v.xunit11-24.vtemp2#branch
.save   v.xunit11-25.vtemp2#branch
.save   v.xunit11-26.vtemp2#branch
.save   v.xunit11-27.vtemp2#branch
.save   v.xunit11-28.vtemp2#branch
.save   v.xunit11-29.vtemp2#branch
.save   v.xunit11-30.vtemp2#branch
.save   v.xunit11-31.vtemp2#branch
.save   v.xunit11-32.vtemp2#branch
.save   v.xunit11-33.vtemp2#branch
.save   v.xunit11-34.vtemp2#branch
.save   v.xunit11-35.vtemp2#branch
.save   v.xunit11-36.vtemp2#branch
.save   v.xunit11-37.vtemp2#branch
.save   v.xunit11-38.vtemp2#branch
.save   v.xunit11-39.vtemp2#branch
.save   v.xunit11-40.vtemp2#branch
.save   v.xunit11-41.vtemp2#branch
.save   v.xunit11-42.vtemp2#branch
.save   v.xunit11-43.vtemp2#branch
.save   v.xunit11-44.vtemp2#branch
.save   v.xunit11-45.vtemp2#branch
.save   v.xunit11-46.vtemp2#branch
.save   v.xunit11-47.vtemp2#branch
.save   v.xunit11-48.vtemp2#branch
.save   v.xunit11-49.vtemp2#branch
.save   v.xunit11-50.vtemp2#branch

.save   v.xunit12-1.vtemp2#branch
.save   v.xunit12-2.vtemp2#branch
.save   v.xunit12-3.vtemp2#branch
.save   v.xunit12-4.vtemp2#branch
.save   v.xunit12-5.vtemp2#branch
.save   v.xunit12-6.vtemp2#branch
.save   v.xunit12-7.vtemp2#branch
.save   v.xunit12-8.vtemp2#branch
.save   v.xunit12-9.vtemp2#branch
.save   v.xunit12-10.vtemp2#branch
.save   v.xunit12-11.vtemp2#branch
.save   v.xunit12-12.vtemp2#branch
.save   v.xunit12-13.vtemp2#branch
.save   v.xunit12-14.vtemp2#branch
.save   v.xunit12-15.vtemp2#branch
.save   v.xunit12-16.vtemp2#branch
.save   v.xunit12-17.vtemp2#branch
.save   v.xunit12-18.vtemp2#branch
.save   v.xunit12-19.vtemp2#branch
.save   v.xunit12-20.vtemp2#branch
.save   v.xunit12-21.vtemp2#branch
.save   v.xunit12-22.vtemp2#branch
.save   v.xunit12-23.vtemp2#branch
.save   v.xunit12-24.vtemp2#branch
.save   v.xunit12-25.vtemp2#branch
.save   v.xunit12-26.vtemp2#branch
.save   v.xunit12-27.vtemp2#branch
.save   v.xunit12-28.vtemp2#branch
.save   v.xunit12-29.vtemp2#branch
.save   v.xunit12-30.vtemp2#branch
.save   v.xunit12-31.vtemp2#branch
.save   v.xunit12-32.vtemp2#branch
.save   v.xunit12-33.vtemp2#branch
.save   v.xunit12-34.vtemp2#branch
.save   v.xunit12-35.vtemp2#branch
.save   v.xunit12-36.vtemp2#branch
.save   v.xunit12-37.vtemp2#branch
.save   v.xunit12-38.vtemp2#branch
.save   v.xunit12-39.vtemp2#branch
.save   v.xunit12-40.vtemp2#branch
.save   v.xunit12-41.vtemp2#branch
.save   v.xunit12-42.vtemp2#branch
.save   v.xunit12-43.vtemp2#branch
.save   v.xunit12-44.vtemp2#branch
.save   v.xunit12-45.vtemp2#branch
.save   v.xunit12-46.vtemp2#branch
.save   v.xunit12-47.vtemp2#branch
.save   v.xunit12-48.vtemp2#branch
.save   v.xunit12-49.vtemp2#branch
.save   v.xunit12-50.vtemp2#branch

.save   v.xunit13-1.vtemp2#branch
.save   v.xunit13-2.vtemp2#branch
.save   v.xunit13-3.vtemp2#branch
.save   v.xunit13-4.vtemp2#branch
.save   v.xunit13-5.vtemp2#branch
.save   v.xunit13-6.vtemp2#branch
.save   v.xunit13-7.vtemp2#branch
.save   v.xunit13-8.vtemp2#branch
.save   v.xunit13-9.vtemp2#branch
.save   v.xunit13-10.vtemp2#branch
.save   v.xunit13-11.vtemp2#branch
.save   v.xunit13-12.vtemp2#branch
.save   v.xunit13-13.vtemp2#branch
.save   v.xunit13-14.vtemp2#branch
.save   v.xunit13-15.vtemp2#branch
.save   v.xunit13-16.vtemp2#branch
.save   v.xunit13-17.vtemp2#branch
.save   v.xunit13-18.vtemp2#branch
.save   v.xunit13-19.vtemp2#branch
.save   v.xunit13-20.vtemp2#branch
.save   v.xunit13-21.vtemp2#branch
.save   v.xunit13-22.vtemp2#branch
.save   v.xunit13-23.vtemp2#branch
.save   v.xunit13-24.vtemp2#branch
.save   v.xunit13-25.vtemp2#branch
.save   v.xunit13-26.vtemp2#branch
.save   v.xunit13-27.vtemp2#branch
.save   v.xunit13-28.vtemp2#branch
.save   v.xunit13-29.vtemp2#branch
.save   v.xunit13-30.vtemp2#branch
.save   v.xunit13-31.vtemp2#branch
.save   v.xunit13-32.vtemp2#branch
.save   v.xunit13-33.vtemp2#branch
.save   v.xunit13-34.vtemp2#branch
.save   v.xunit13-35.vtemp2#branch
.save   v.xunit13-36.vtemp2#branch
.save   v.xunit13-37.vtemp2#branch
.save   v.xunit13-38.vtemp2#branch
.save   v.xunit13-39.vtemp2#branch
.save   v.xunit13-40.vtemp2#branch
.save   v.xunit13-41.vtemp2#branch
.save   v.xunit13-42.vtemp2#branch
.save   v.xunit13-43.vtemp2#branch
.save   v.xunit13-44.vtemp2#branch
.save   v.xunit13-45.vtemp2#branch
.save   v.xunit13-46.vtemp2#branch
.save   v.xunit13-47.vtemp2#branch
.save   v.xunit13-48.vtemp2#branch
.save   v.xunit13-49.vtemp2#branch
.save   v.xunit13-50.vtemp2#branch

.save   v.xunit14-1.vtemp2#branch
.save   v.xunit14-2.vtemp2#branch
.save   v.xunit14-3.vtemp2#branch
.save   v.xunit14-4.vtemp2#branch
.save   v.xunit14-5.vtemp2#branch
.save   v.xunit14-6.vtemp2#branch
.save   v.xunit14-7.vtemp2#branch
.save   v.xunit14-8.vtemp2#branch
.save   v.xunit14-9.vtemp2#branch
.save   v.xunit14-10.vtemp2#branch
.save   v.xunit14-11.vtemp2#branch
.save   v.xunit14-12.vtemp2#branch
.save   v.xunit14-13.vtemp2#branch
.save   v.xunit14-14.vtemp2#branch
.save   v.xunit14-15.vtemp2#branch
.save   v.xunit14-16.vtemp2#branch
.save   v.xunit14-17.vtemp2#branch
.save   v.xunit14-18.vtemp2#branch
.save   v.xunit14-19.vtemp2#branch
.save   v.xunit14-20.vtemp2#branch
.save   v.xunit14-21.vtemp2#branch
.save   v.xunit14-22.vtemp2#branch
.save   v.xunit14-23.vtemp2#branch
.save   v.xunit14-24.vtemp2#branch
.save   v.xunit14-25.vtemp2#branch
.save   v.xunit14-26.vtemp2#branch
.save   v.xunit14-27.vtemp2#branch
.save   v.xunit14-28.vtemp2#branch
.save   v.xunit14-29.vtemp2#branch
.save   v.xunit14-30.vtemp2#branch
.save   v.xunit14-31.vtemp2#branch
.save   v.xunit14-32.vtemp2#branch
.save   v.xunit14-33.vtemp2#branch
.save   v.xunit14-34.vtemp2#branch
.save   v.xunit14-35.vtemp2#branch
.save   v.xunit14-36.vtemp2#branch
.save   v.xunit14-37.vtemp2#branch
.save   v.xunit14-38.vtemp2#branch
.save   v.xunit14-39.vtemp2#branch
.save   v.xunit14-40.vtemp2#branch
.save   v.xunit14-41.vtemp2#branch
.save   v.xunit14-42.vtemp2#branch
.save   v.xunit14-43.vtemp2#branch
.save   v.xunit14-44.vtemp2#branch
.save   v.xunit14-45.vtemp2#branch
.save   v.xunit14-46.vtemp2#branch
.save   v.xunit14-47.vtemp2#branch
.save   v.xunit14-48.vtemp2#branch
.save   v.xunit14-49.vtemp2#branch
.save   v.xunit14-50.vtemp2#branch

.save   v.xunit15-1.vtemp2#branch
.save   v.xunit15-2.vtemp2#branch
.save   v.xunit15-3.vtemp2#branch
.save   v.xunit15-4.vtemp2#branch
.save   v.xunit15-5.vtemp2#branch
.save   v.xunit15-6.vtemp2#branch
.save   v.xunit15-7.vtemp2#branch
.save   v.xunit15-8.vtemp2#branch
.save   v.xunit15-9.vtemp2#branch
.save   v.xunit15-10.vtemp2#branch
.save   v.xunit15-11.vtemp2#branch
.save   v.xunit15-12.vtemp2#branch
.save   v.xunit15-13.vtemp2#branch
.save   v.xunit15-14.vtemp2#branch
.save   v.xunit15-15.vtemp2#branch
.save   v.xunit15-16.vtemp2#branch
.save   v.xunit15-17.vtemp2#branch
.save   v.xunit15-18.vtemp2#branch
.save   v.xunit15-19.vtemp2#branch
.save   v.xunit15-20.vtemp2#branch
.save   v.xunit15-21.vtemp2#branch
.save   v.xunit15-22.vtemp2#branch
.save   v.xunit15-23.vtemp2#branch
.save   v.xunit15-24.vtemp2#branch
.save   v.xunit15-25.vtemp2#branch
.save   v.xunit15-26.vtemp2#branch
.save   v.xunit15-27.vtemp2#branch
.save   v.xunit15-28.vtemp2#branch
.save   v.xunit15-29.vtemp2#branch
.save   v.xunit15-30.vtemp2#branch
.save   v.xunit15-31.vtemp2#branch
.save   v.xunit15-32.vtemp2#branch
.save   v.xunit15-33.vtemp2#branch
.save   v.xunit15-34.vtemp2#branch
.save   v.xunit15-35.vtemp2#branch
.save   v.xunit15-36.vtemp2#branch
.save   v.xunit15-37.vtemp2#branch
.save   v.xunit15-38.vtemp2#branch
.save   v.xunit15-39.vtemp2#branch
.save   v.xunit15-40.vtemp2#branch
.save   v.xunit15-41.vtemp2#branch
.save   v.xunit15-42.vtemp2#branch
.save   v.xunit15-43.vtemp2#branch
.save   v.xunit15-44.vtemp2#branch
.save   v.xunit15-45.vtemp2#branch
.save   v.xunit15-46.vtemp2#branch
.save   v.xunit15-47.vtemp2#branch
.save   v.xunit15-48.vtemp2#branch
.save   v.xunit15-49.vtemp2#branch
.save   v.xunit15-50.vtemp2#branch

.save   v.xunit16-1.vtemp2#branch
.save   v.xunit16-2.vtemp2#branch
.save   v.xunit16-3.vtemp2#branch
.save   v.xunit16-4.vtemp2#branch
.save   v.xunit16-5.vtemp2#branch
.save   v.xunit16-6.vtemp2#branch
.save   v.xunit16-7.vtemp2#branch
.save   v.xunit16-8.vtemp2#branch
.save   v.xunit16-9.vtemp2#branch
.save   v.xunit16-10.vtemp2#branch
.save   v.xunit16-11.vtemp2#branch
.save   v.xunit16-12.vtemp2#branch
.save   v.xunit16-13.vtemp2#branch
.save   v.xunit16-14.vtemp2#branch
.save   v.xunit16-15.vtemp2#branch
.save   v.xunit16-16.vtemp2#branch
.save   v.xunit16-17.vtemp2#branch
.save   v.xunit16-18.vtemp2#branch
.save   v.xunit16-19.vtemp2#branch
.save   v.xunit16-20.vtemp2#branch
.save   v.xunit16-21.vtemp2#branch
.save   v.xunit16-22.vtemp2#branch
.save   v.xunit16-23.vtemp2#branch
.save   v.xunit16-24.vtemp2#branch
.save   v.xunit16-25.vtemp2#branch
.save   v.xunit16-26.vtemp2#branch
.save   v.xunit16-27.vtemp2#branch
.save   v.xunit16-28.vtemp2#branch
.save   v.xunit16-29.vtemp2#branch
.save   v.xunit16-30.vtemp2#branch
.save   v.xunit16-31.vtemp2#branch
.save   v.xunit16-32.vtemp2#branch
.save   v.xunit16-33.vtemp2#branch
.save   v.xunit16-34.vtemp2#branch
.save   v.xunit16-35.vtemp2#branch
.save   v.xunit16-36.vtemp2#branch
.save   v.xunit16-37.vtemp2#branch
.save   v.xunit16-38.vtemp2#branch
.save   v.xunit16-39.vtemp2#branch
.save   v.xunit16-40.vtemp2#branch
.save   v.xunit16-41.vtemp2#branch
.save   v.xunit16-42.vtemp2#branch
.save   v.xunit16-43.vtemp2#branch
.save   v.xunit16-44.vtemp2#branch
.save   v.xunit16-45.vtemp2#branch
.save   v.xunit16-46.vtemp2#branch
.save   v.xunit16-47.vtemp2#branch
.save   v.xunit16-48.vtemp2#branch
.save   v.xunit16-49.vtemp2#branch
.save   v.xunit16-50.vtemp2#branch

.save   v.xunit17-1.vtemp2#branch
.save   v.xunit17-2.vtemp2#branch
.save   v.xunit17-3.vtemp2#branch
.save   v.xunit17-4.vtemp2#branch
.save   v.xunit17-5.vtemp2#branch
.save   v.xunit17-6.vtemp2#branch
.save   v.xunit17-7.vtemp2#branch
.save   v.xunit17-8.vtemp2#branch
.save   v.xunit17-9.vtemp2#branch
.save   v.xunit17-10.vtemp2#branch
.save   v.xunit17-11.vtemp2#branch
.save   v.xunit17-12.vtemp2#branch
.save   v.xunit17-13.vtemp2#branch
.save   v.xunit17-14.vtemp2#branch
.save   v.xunit17-15.vtemp2#branch
.save   v.xunit17-16.vtemp2#branch
.save   v.xunit17-17.vtemp2#branch
.save   v.xunit17-18.vtemp2#branch
.save   v.xunit17-19.vtemp2#branch
.save   v.xunit17-20.vtemp2#branch
.save   v.xunit17-21.vtemp2#branch
.save   v.xunit17-22.vtemp2#branch
.save   v.xunit17-23.vtemp2#branch
.save   v.xunit17-24.vtemp2#branch
.save   v.xunit17-25.vtemp2#branch
.save   v.xunit17-26.vtemp2#branch
.save   v.xunit17-27.vtemp2#branch
.save   v.xunit17-28.vtemp2#branch
.save   v.xunit17-29.vtemp2#branch
.save   v.xunit17-30.vtemp2#branch
.save   v.xunit17-31.vtemp2#branch
.save   v.xunit17-32.vtemp2#branch
.save   v.xunit17-33.vtemp2#branch
.save   v.xunit17-34.vtemp2#branch
.save   v.xunit17-35.vtemp2#branch
.save   v.xunit17-36.vtemp2#branch
.save   v.xunit17-37.vtemp2#branch
.save   v.xunit17-38.vtemp2#branch
.save   v.xunit17-39.vtemp2#branch
.save   v.xunit17-40.vtemp2#branch
.save   v.xunit17-41.vtemp2#branch
.save   v.xunit17-42.vtemp2#branch
.save   v.xunit17-43.vtemp2#branch
.save   v.xunit17-44.vtemp2#branch
.save   v.xunit17-45.vtemp2#branch
.save   v.xunit17-46.vtemp2#branch
.save   v.xunit17-47.vtemp2#branch
.save   v.xunit17-48.vtemp2#branch
.save   v.xunit17-49.vtemp2#branch
.save   v.xunit17-50.vtemp2#branch

.save   v.xunit18-1.vtemp2#branch
.save   v.xunit18-2.vtemp2#branch
.save   v.xunit18-3.vtemp2#branch
.save   v.xunit18-4.vtemp2#branch
.save   v.xunit18-5.vtemp2#branch
.save   v.xunit18-6.vtemp2#branch
.save   v.xunit18-7.vtemp2#branch
.save   v.xunit18-8.vtemp2#branch
.save   v.xunit18-9.vtemp2#branch
.save   v.xunit18-10.vtemp2#branch
.save   v.xunit18-11.vtemp2#branch
.save   v.xunit18-12.vtemp2#branch
.save   v.xunit18-13.vtemp2#branch
.save   v.xunit18-14.vtemp2#branch
.save   v.xunit18-15.vtemp2#branch
.save   v.xunit18-16.vtemp2#branch
.save   v.xunit18-17.vtemp2#branch
.save   v.xunit18-18.vtemp2#branch
.save   v.xunit18-19.vtemp2#branch
.save   v.xunit18-20.vtemp2#branch
.save   v.xunit18-21.vtemp2#branch
.save   v.xunit18-22.vtemp2#branch
.save   v.xunit18-23.vtemp2#branch
.save   v.xunit18-24.vtemp2#branch
.save   v.xunit18-25.vtemp2#branch
.save   v.xunit18-26.vtemp2#branch
.save   v.xunit18-27.vtemp2#branch
.save   v.xunit18-28.vtemp2#branch
.save   v.xunit18-29.vtemp2#branch
.save   v.xunit18-30.vtemp2#branch
.save   v.xunit18-31.vtemp2#branch
.save   v.xunit18-32.vtemp2#branch
.save   v.xunit18-33.vtemp2#branch
.save   v.xunit18-34.vtemp2#branch
.save   v.xunit18-35.vtemp2#branch
.save   v.xunit18-36.vtemp2#branch
.save   v.xunit18-37.vtemp2#branch
.save   v.xunit18-38.vtemp2#branch
.save   v.xunit18-39.vtemp2#branch
.save   v.xunit18-40.vtemp2#branch
.save   v.xunit18-41.vtemp2#branch
.save   v.xunit18-42.vtemp2#branch
.save   v.xunit18-43.vtemp2#branch
.save   v.xunit18-44.vtemp2#branch
.save   v.xunit18-45.vtemp2#branch
.save   v.xunit18-46.vtemp2#branch
.save   v.xunit18-47.vtemp2#branch
.save   v.xunit18-48.vtemp2#branch
.save   v.xunit18-49.vtemp2#branch
.save   v.xunit18-50.vtemp2#branch

.save   v.xunit19-1.vtemp2#branch
.save   v.xunit19-2.vtemp2#branch
.save   v.xunit19-3.vtemp2#branch
.save   v.xunit19-4.vtemp2#branch
.save   v.xunit19-5.vtemp2#branch
.save   v.xunit19-6.vtemp2#branch
.save   v.xunit19-7.vtemp2#branch
.save   v.xunit19-8.vtemp2#branch
.save   v.xunit19-9.vtemp2#branch
.save   v.xunit19-10.vtemp2#branch
.save   v.xunit19-11.vtemp2#branch
.save   v.xunit19-12.vtemp2#branch
.save   v.xunit19-13.vtemp2#branch
.save   v.xunit19-14.vtemp2#branch
.save   v.xunit19-15.vtemp2#branch
.save   v.xunit19-16.vtemp2#branch
.save   v.xunit19-17.vtemp2#branch
.save   v.xunit19-18.vtemp2#branch
.save   v.xunit19-19.vtemp2#branch
.save   v.xunit19-20.vtemp2#branch
.save   v.xunit19-21.vtemp2#branch
.save   v.xunit19-22.vtemp2#branch
.save   v.xunit19-23.vtemp2#branch
.save   v.xunit19-24.vtemp2#branch
.save   v.xunit19-25.vtemp2#branch
.save   v.xunit19-26.vtemp2#branch
.save   v.xunit19-27.vtemp2#branch
.save   v.xunit19-28.vtemp2#branch
.save   v.xunit19-29.vtemp2#branch
.save   v.xunit19-30.vtemp2#branch
.save   v.xunit19-31.vtemp2#branch
.save   v.xunit19-32.vtemp2#branch
.save   v.xunit19-33.vtemp2#branch
.save   v.xunit19-34.vtemp2#branch
.save   v.xunit19-35.vtemp2#branch
.save   v.xunit19-36.vtemp2#branch
.save   v.xunit19-37.vtemp2#branch
.save   v.xunit19-38.vtemp2#branch
.save   v.xunit19-39.vtemp2#branch
.save   v.xunit19-40.vtemp2#branch
.save   v.xunit19-41.vtemp2#branch
.save   v.xunit19-42.vtemp2#branch
.save   v.xunit19-43.vtemp2#branch
.save   v.xunit19-44.vtemp2#branch
.save   v.xunit19-45.vtemp2#branch
.save   v.xunit19-46.vtemp2#branch
.save   v.xunit19-47.vtemp2#branch
.save   v.xunit19-48.vtemp2#branch
.save   v.xunit19-49.vtemp2#branch
.save   v.xunit19-50.vtemp2#branch

.save   v.xunit20-1.vtemp2#branch
.save   v.xunit20-2.vtemp2#branch
.save   v.xunit20-3.vtemp2#branch
.save   v.xunit20-4.vtemp2#branch
.save   v.xunit20-5.vtemp2#branch
.save   v.xunit20-6.vtemp2#branch
.save   v.xunit20-7.vtemp2#branch
.save   v.xunit20-8.vtemp2#branch
.save   v.xunit20-9.vtemp2#branch
.save   v.xunit20-10.vtemp2#branch
.save   v.xunit20-11.vtemp2#branch
.save   v.xunit20-12.vtemp2#branch
.save   v.xunit20-13.vtemp2#branch
.save   v.xunit20-14.vtemp2#branch
.save   v.xunit20-15.vtemp2#branch
.save   v.xunit20-16.vtemp2#branch
.save   v.xunit20-17.vtemp2#branch
.save   v.xunit20-18.vtemp2#branch
.save   v.xunit20-19.vtemp2#branch
.save   v.xunit20-20.vtemp2#branch
.save   v.xunit20-21.vtemp2#branch
.save   v.xunit20-22.vtemp2#branch
.save   v.xunit20-23.vtemp2#branch
.save   v.xunit20-24.vtemp2#branch
.save   v.xunit20-25.vtemp2#branch
.save   v.xunit20-26.vtemp2#branch
.save   v.xunit20-27.vtemp2#branch
.save   v.xunit20-28.vtemp2#branch
.save   v.xunit20-29.vtemp2#branch
.save   v.xunit20-30.vtemp2#branch
.save   v.xunit20-31.vtemp2#branch
.save   v.xunit20-32.vtemp2#branch
.save   v.xunit20-33.vtemp2#branch
.save   v.xunit20-34.vtemp2#branch
.save   v.xunit20-35.vtemp2#branch
.save   v.xunit20-36.vtemp2#branch
.save   v.xunit20-37.vtemp2#branch
.save   v.xunit20-38.vtemp2#branch
.save   v.xunit20-39.vtemp2#branch
.save   v.xunit20-40.vtemp2#branch
.save   v.xunit20-41.vtemp2#branch
.save   v.xunit20-42.vtemp2#branch
.save   v.xunit20-43.vtemp2#branch
.save   v.xunit20-44.vtemp2#branch
.save   v.xunit20-45.vtemp2#branch
.save   v.xunit20-46.vtemp2#branch
.save   v.xunit20-47.vtemp2#branch
.save   v.xunit20-48.vtemp2#branch
.save   v.xunit20-49.vtemp2#branch
.save   v.xunit20-50.vtemp2#branch

.save   v.xunit21-1.vtemp2#branch
.save   v.xunit21-2.vtemp2#branch
.save   v.xunit21-3.vtemp2#branch
.save   v.xunit21-4.vtemp2#branch
.save   v.xunit21-5.vtemp2#branch
.save   v.xunit21-6.vtemp2#branch
.save   v.xunit21-7.vtemp2#branch
.save   v.xunit21-8.vtemp2#branch
.save   v.xunit21-9.vtemp2#branch
.save   v.xunit21-10.vtemp2#branch
.save   v.xunit21-11.vtemp2#branch
.save   v.xunit21-12.vtemp2#branch
.save   v.xunit21-13.vtemp2#branch
.save   v.xunit21-14.vtemp2#branch
.save   v.xunit21-15.vtemp2#branch
.save   v.xunit21-16.vtemp2#branch
.save   v.xunit21-17.vtemp2#branch
.save   v.xunit21-18.vtemp2#branch
.save   v.xunit21-19.vtemp2#branch
.save   v.xunit21-20.vtemp2#branch
.save   v.xunit21-21.vtemp2#branch
.save   v.xunit21-22.vtemp2#branch
.save   v.xunit21-23.vtemp2#branch
.save   v.xunit21-24.vtemp2#branch
.save   v.xunit21-25.vtemp2#branch
.save   v.xunit21-26.vtemp2#branch
.save   v.xunit21-27.vtemp2#branch
.save   v.xunit21-28.vtemp2#branch
.save   v.xunit21-29.vtemp2#branch
.save   v.xunit21-30.vtemp2#branch
.save   v.xunit21-31.vtemp2#branch
.save   v.xunit21-32.vtemp2#branch
.save   v.xunit21-33.vtemp2#branch
.save   v.xunit21-34.vtemp2#branch
.save   v.xunit21-35.vtemp2#branch
.save   v.xunit21-36.vtemp2#branch
.save   v.xunit21-37.vtemp2#branch
.save   v.xunit21-38.vtemp2#branch
.save   v.xunit21-39.vtemp2#branch
.save   v.xunit21-40.vtemp2#branch
.save   v.xunit21-41.vtemp2#branch
.save   v.xunit21-42.vtemp2#branch
.save   v.xunit21-43.vtemp2#branch
.save   v.xunit21-44.vtemp2#branch
.save   v.xunit21-45.vtemp2#branch
.save   v.xunit21-46.vtemp2#branch
.save   v.xunit21-47.vtemp2#branch
.save   v.xunit21-48.vtemp2#branch
.save   v.xunit21-49.vtemp2#branch
.save   v.xunit21-50.vtemp2#branch

.save   v.xunit22-1.vtemp2#branch
.save   v.xunit22-2.vtemp2#branch
.save   v.xunit22-3.vtemp2#branch
.save   v.xunit22-4.vtemp2#branch
.save   v.xunit22-5.vtemp2#branch
.save   v.xunit22-6.vtemp2#branch
.save   v.xunit22-7.vtemp2#branch
.save   v.xunit22-8.vtemp2#branch
.save   v.xunit22-9.vtemp2#branch
.save   v.xunit22-10.vtemp2#branch
.save   v.xunit22-11.vtemp2#branch
.save   v.xunit22-12.vtemp2#branch
.save   v.xunit22-13.vtemp2#branch
.save   v.xunit22-14.vtemp2#branch
.save   v.xunit22-15.vtemp2#branch
.save   v.xunit22-16.vtemp2#branch
.save   v.xunit22-17.vtemp2#branch
.save   v.xunit22-18.vtemp2#branch
.save   v.xunit22-19.vtemp2#branch
.save   v.xunit22-20.vtemp2#branch
.save   v.xunit22-21.vtemp2#branch
.save   v.xunit22-22.vtemp2#branch
.save   v.xunit22-23.vtemp2#branch
.save   v.xunit22-24.vtemp2#branch
.save   v.xunit22-25.vtemp2#branch
.save   v.xunit22-26.vtemp2#branch
.save   v.xunit22-27.vtemp2#branch
.save   v.xunit22-28.vtemp2#branch
.save   v.xunit22-29.vtemp2#branch
.save   v.xunit22-30.vtemp2#branch
.save   v.xunit22-31.vtemp2#branch
.save   v.xunit22-32.vtemp2#branch
.save   v.xunit22-33.vtemp2#branch
.save   v.xunit22-34.vtemp2#branch
.save   v.xunit22-35.vtemp2#branch
.save   v.xunit22-36.vtemp2#branch
.save   v.xunit22-37.vtemp2#branch
.save   v.xunit22-38.vtemp2#branch
.save   v.xunit22-39.vtemp2#branch
.save   v.xunit22-40.vtemp2#branch
.save   v.xunit22-41.vtemp2#branch
.save   v.xunit22-42.vtemp2#branch
.save   v.xunit22-43.vtemp2#branch
.save   v.xunit22-44.vtemp2#branch
.save   v.xunit22-45.vtemp2#branch
.save   v.xunit22-46.vtemp2#branch
.save   v.xunit22-47.vtemp2#branch
.save   v.xunit22-48.vtemp2#branch
.save   v.xunit22-49.vtemp2#branch
.save   v.xunit22-50.vtemp2#branch

.save   v.xunit23-1.vtemp2#branch
.save   v.xunit23-2.vtemp2#branch
.save   v.xunit23-3.vtemp2#branch
.save   v.xunit23-4.vtemp2#branch
.save   v.xunit23-5.vtemp2#branch
.save   v.xunit23-6.vtemp2#branch
.save   v.xunit23-7.vtemp2#branch
.save   v.xunit23-8.vtemp2#branch
.save   v.xunit23-9.vtemp2#branch
.save   v.xunit23-10.vtemp2#branch
.save   v.xunit23-11.vtemp2#branch
.save   v.xunit23-12.vtemp2#branch
.save   v.xunit23-13.vtemp2#branch
.save   v.xunit23-14.vtemp2#branch
.save   v.xunit23-15.vtemp2#branch
.save   v.xunit23-16.vtemp2#branch
.save   v.xunit23-17.vtemp2#branch
.save   v.xunit23-18.vtemp2#branch
.save   v.xunit23-19.vtemp2#branch
.save   v.xunit23-20.vtemp2#branch
.save   v.xunit23-21.vtemp2#branch
.save   v.xunit23-22.vtemp2#branch
.save   v.xunit23-23.vtemp2#branch
.save   v.xunit23-24.vtemp2#branch
.save   v.xunit23-25.vtemp2#branch
.save   v.xunit23-26.vtemp2#branch
.save   v.xunit23-27.vtemp2#branch
.save   v.xunit23-28.vtemp2#branch
.save   v.xunit23-29.vtemp2#branch
.save   v.xunit23-30.vtemp2#branch
.save   v.xunit23-31.vtemp2#branch
.save   v.xunit23-32.vtemp2#branch
.save   v.xunit23-33.vtemp2#branch
.save   v.xunit23-34.vtemp2#branch
.save   v.xunit23-35.vtemp2#branch
.save   v.xunit23-36.vtemp2#branch
.save   v.xunit23-37.vtemp2#branch
.save   v.xunit23-38.vtemp2#branch
.save   v.xunit23-39.vtemp2#branch
.save   v.xunit23-40.vtemp2#branch
.save   v.xunit23-41.vtemp2#branch
.save   v.xunit23-42.vtemp2#branch
.save   v.xunit23-43.vtemp2#branch
.save   v.xunit23-44.vtemp2#branch
.save   v.xunit23-45.vtemp2#branch
.save   v.xunit23-46.vtemp2#branch
.save   v.xunit23-47.vtemp2#branch
.save   v.xunit23-48.vtemp2#branch
.save   v.xunit23-49.vtemp2#branch
.save   v.xunit23-50.vtemp2#branch

.save   v.xunit24-1.vtemp2#branch
.save   v.xunit24-2.vtemp2#branch
.save   v.xunit24-3.vtemp2#branch
.save   v.xunit24-4.vtemp2#branch
.save   v.xunit24-5.vtemp2#branch
.save   v.xunit24-6.vtemp2#branch
.save   v.xunit24-7.vtemp2#branch
.save   v.xunit24-8.vtemp2#branch
.save   v.xunit24-9.vtemp2#branch
.save   v.xunit24-10.vtemp2#branch
.save   v.xunit24-11.vtemp2#branch
.save   v.xunit24-12.vtemp2#branch
.save   v.xunit24-13.vtemp2#branch
.save   v.xunit24-14.vtemp2#branch
.save   v.xunit24-15.vtemp2#branch
.save   v.xunit24-16.vtemp2#branch
.save   v.xunit24-17.vtemp2#branch
.save   v.xunit24-18.vtemp2#branch
.save   v.xunit24-19.vtemp2#branch
.save   v.xunit24-20.vtemp2#branch
.save   v.xunit24-21.vtemp2#branch
.save   v.xunit24-22.vtemp2#branch
.save   v.xunit24-23.vtemp2#branch
.save   v.xunit24-24.vtemp2#branch
.save   v.xunit24-25.vtemp2#branch
.save   v.xunit24-26.vtemp2#branch
.save   v.xunit24-27.vtemp2#branch
.save   v.xunit24-28.vtemp2#branch
.save   v.xunit24-29.vtemp2#branch
.save   v.xunit24-30.vtemp2#branch
.save   v.xunit24-31.vtemp2#branch
.save   v.xunit24-32.vtemp2#branch
.save   v.xunit24-33.vtemp2#branch
.save   v.xunit24-34.vtemp2#branch
.save   v.xunit24-35.vtemp2#branch
.save   v.xunit24-36.vtemp2#branch
.save   v.xunit24-37.vtemp2#branch
.save   v.xunit24-38.vtemp2#branch
.save   v.xunit24-39.vtemp2#branch
.save   v.xunit24-40.vtemp2#branch
.save   v.xunit24-41.vtemp2#branch
.save   v.xunit24-42.vtemp2#branch
.save   v.xunit24-43.vtemp2#branch
.save   v.xunit24-44.vtemp2#branch
.save   v.xunit24-45.vtemp2#branch
.save   v.xunit24-46.vtemp2#branch
.save   v.xunit24-47.vtemp2#branch
.save   v.xunit24-48.vtemp2#branch
.save   v.xunit24-49.vtemp2#branch
.save   v.xunit24-50.vtemp2#branch

.save   v.xunit25-1.vtemp2#branch
.save   v.xunit25-2.vtemp2#branch
.save   v.xunit25-3.vtemp2#branch
.save   v.xunit25-4.vtemp2#branch
.save   v.xunit25-5.vtemp2#branch
.save   v.xunit25-6.vtemp2#branch
.save   v.xunit25-7.vtemp2#branch
.save   v.xunit25-8.vtemp2#branch
.save   v.xunit25-9.vtemp2#branch
.save   v.xunit25-10.vtemp2#branch
.save   v.xunit25-11.vtemp2#branch
.save   v.xunit25-12.vtemp2#branch
.save   v.xunit25-13.vtemp2#branch
.save   v.xunit25-14.vtemp2#branch
.save   v.xunit25-15.vtemp2#branch
.save   v.xunit25-16.vtemp2#branch
.save   v.xunit25-17.vtemp2#branch
.save   v.xunit25-18.vtemp2#branch
.save   v.xunit25-19.vtemp2#branch
.save   v.xunit25-20.vtemp2#branch
.save   v.xunit25-21.vtemp2#branch
.save   v.xunit25-22.vtemp2#branch
.save   v.xunit25-23.vtemp2#branch
.save   v.xunit25-24.vtemp2#branch
.save   v.xunit25-25.vtemp2#branch
.save   v.xunit25-26.vtemp2#branch
.save   v.xunit25-27.vtemp2#branch
.save   v.xunit25-28.vtemp2#branch
.save   v.xunit25-29.vtemp2#branch
.save   v.xunit25-30.vtemp2#branch
.save   v.xunit25-31.vtemp2#branch
.save   v.xunit25-32.vtemp2#branch
.save   v.xunit25-33.vtemp2#branch
.save   v.xunit25-34.vtemp2#branch
.save   v.xunit25-35.vtemp2#branch
.save   v.xunit25-36.vtemp2#branch
.save   v.xunit25-37.vtemp2#branch
.save   v.xunit25-38.vtemp2#branch
.save   v.xunit25-39.vtemp2#branch
.save   v.xunit25-40.vtemp2#branch
.save   v.xunit25-41.vtemp2#branch
.save   v.xunit25-42.vtemp2#branch
.save   v.xunit25-43.vtemp2#branch
.save   v.xunit25-44.vtemp2#branch
.save   v.xunit25-45.vtemp2#branch
.save   v.xunit25-46.vtemp2#branch
.save   v.xunit25-47.vtemp2#branch
.save   v.xunit25-48.vtemp2#branch
.save   v.xunit25-49.vtemp2#branch
.save   v.xunit25-50.vtemp2#branch

.save   v.xunit26-1.vtemp2#branch
.save   v.xunit26-2.vtemp2#branch
.save   v.xunit26-3.vtemp2#branch
.save   v.xunit26-4.vtemp2#branch
.save   v.xunit26-5.vtemp2#branch
.save   v.xunit26-6.vtemp2#branch
.save   v.xunit26-7.vtemp2#branch
.save   v.xunit26-8.vtemp2#branch
.save   v.xunit26-9.vtemp2#branch
.save   v.xunit26-10.vtemp2#branch
.save   v.xunit26-11.vtemp2#branch
.save   v.xunit26-12.vtemp2#branch
.save   v.xunit26-13.vtemp2#branch
.save   v.xunit26-14.vtemp2#branch
.save   v.xunit26-15.vtemp2#branch
.save   v.xunit26-16.vtemp2#branch
.save   v.xunit26-17.vtemp2#branch
.save   v.xunit26-18.vtemp2#branch
.save   v.xunit26-19.vtemp2#branch
.save   v.xunit26-20.vtemp2#branch
.save   v.xunit26-21.vtemp2#branch
.save   v.xunit26-22.vtemp2#branch
.save   v.xunit26-23.vtemp2#branch
.save   v.xunit26-24.vtemp2#branch
.save   v.xunit26-25.vtemp2#branch
.save   v.xunit26-26.vtemp2#branch
.save   v.xunit26-27.vtemp2#branch
.save   v.xunit26-28.vtemp2#branch
.save   v.xunit26-29.vtemp2#branch
.save   v.xunit26-30.vtemp2#branch
.save   v.xunit26-31.vtemp2#branch
.save   v.xunit26-32.vtemp2#branch
.save   v.xunit26-33.vtemp2#branch
.save   v.xunit26-34.vtemp2#branch
.save   v.xunit26-35.vtemp2#branch
.save   v.xunit26-36.vtemp2#branch
.save   v.xunit26-37.vtemp2#branch
.save   v.xunit26-38.vtemp2#branch
.save   v.xunit26-39.vtemp2#branch
.save   v.xunit26-40.vtemp2#branch
.save   v.xunit26-41.vtemp2#branch
.save   v.xunit26-42.vtemp2#branch
.save   v.xunit26-43.vtemp2#branch
.save   v.xunit26-44.vtemp2#branch
.save   v.xunit26-45.vtemp2#branch
.save   v.xunit26-46.vtemp2#branch
.save   v.xunit26-47.vtemp2#branch
.save   v.xunit26-48.vtemp2#branch
.save   v.xunit26-49.vtemp2#branch
.save   v.xunit26-50.vtemp2#branch

.save   v.xunit27-1.vtemp2#branch
.save   v.xunit27-2.vtemp2#branch
.save   v.xunit27-3.vtemp2#branch
.save   v.xunit27-4.vtemp2#branch
.save   v.xunit27-5.vtemp2#branch
.save   v.xunit27-6.vtemp2#branch
.save   v.xunit27-7.vtemp2#branch
.save   v.xunit27-8.vtemp2#branch
.save   v.xunit27-9.vtemp2#branch
.save   v.xunit27-10.vtemp2#branch
.save   v.xunit27-11.vtemp2#branch
.save   v.xunit27-12.vtemp2#branch
.save   v.xunit27-13.vtemp2#branch
.save   v.xunit27-14.vtemp2#branch
.save   v.xunit27-15.vtemp2#branch
.save   v.xunit27-16.vtemp2#branch
.save   v.xunit27-17.vtemp2#branch
.save   v.xunit27-18.vtemp2#branch
.save   v.xunit27-19.vtemp2#branch
.save   v.xunit27-20.vtemp2#branch
.save   v.xunit27-21.vtemp2#branch
.save   v.xunit27-22.vtemp2#branch
.save   v.xunit27-23.vtemp2#branch
.save   v.xunit27-24.vtemp2#branch
.save   v.xunit27-25.vtemp2#branch
.save   v.xunit27-26.vtemp2#branch
.save   v.xunit27-27.vtemp2#branch
.save   v.xunit27-28.vtemp2#branch
.save   v.xunit27-29.vtemp2#branch
.save   v.xunit27-30.vtemp2#branch
.save   v.xunit27-31.vtemp2#branch
.save   v.xunit27-32.vtemp2#branch
.save   v.xunit27-33.vtemp2#branch
.save   v.xunit27-34.vtemp2#branch
.save   v.xunit27-35.vtemp2#branch
.save   v.xunit27-36.vtemp2#branch
.save   v.xunit27-37.vtemp2#branch
.save   v.xunit27-38.vtemp2#branch
.save   v.xunit27-39.vtemp2#branch
.save   v.xunit27-40.vtemp2#branch
.save   v.xunit27-41.vtemp2#branch
.save   v.xunit27-42.vtemp2#branch
.save   v.xunit27-43.vtemp2#branch
.save   v.xunit27-44.vtemp2#branch
.save   v.xunit27-45.vtemp2#branch
.save   v.xunit27-46.vtemp2#branch
.save   v.xunit27-47.vtemp2#branch
.save   v.xunit27-48.vtemp2#branch
.save   v.xunit27-49.vtemp2#branch
.save   v.xunit27-50.vtemp2#branch

.save   v.xunit28-1.vtemp2#branch
.save   v.xunit28-2.vtemp2#branch
.save   v.xunit28-3.vtemp2#branch
.save   v.xunit28-4.vtemp2#branch
.save   v.xunit28-5.vtemp2#branch
.save   v.xunit28-6.vtemp2#branch
.save   v.xunit28-7.vtemp2#branch
.save   v.xunit28-8.vtemp2#branch
.save   v.xunit28-9.vtemp2#branch
.save   v.xunit28-10.vtemp2#branch
.save   v.xunit28-11.vtemp2#branch
.save   v.xunit28-12.vtemp2#branch
.save   v.xunit28-13.vtemp2#branch
.save   v.xunit28-14.vtemp2#branch
.save   v.xunit28-15.vtemp2#branch
.save   v.xunit28-16.vtemp2#branch
.save   v.xunit28-17.vtemp2#branch
.save   v.xunit28-18.vtemp2#branch
.save   v.xunit28-19.vtemp2#branch
.save   v.xunit28-20.vtemp2#branch
.save   v.xunit28-21.vtemp2#branch
.save   v.xunit28-22.vtemp2#branch
.save   v.xunit28-23.vtemp2#branch
.save   v.xunit28-24.vtemp2#branch
.save   v.xunit28-25.vtemp2#branch
.save   v.xunit28-26.vtemp2#branch
.save   v.xunit28-27.vtemp2#branch
.save   v.xunit28-28.vtemp2#branch
.save   v.xunit28-29.vtemp2#branch
.save   v.xunit28-30.vtemp2#branch
.save   v.xunit28-31.vtemp2#branch
.save   v.xunit28-32.vtemp2#branch
.save   v.xunit28-33.vtemp2#branch
.save   v.xunit28-34.vtemp2#branch
.save   v.xunit28-35.vtemp2#branch
.save   v.xunit28-36.vtemp2#branch
.save   v.xunit28-37.vtemp2#branch
.save   v.xunit28-38.vtemp2#branch
.save   v.xunit28-39.vtemp2#branch
.save   v.xunit28-40.vtemp2#branch
.save   v.xunit28-41.vtemp2#branch
.save   v.xunit28-42.vtemp2#branch
.save   v.xunit28-43.vtemp2#branch
.save   v.xunit28-44.vtemp2#branch
.save   v.xunit28-45.vtemp2#branch
.save   v.xunit28-46.vtemp2#branch
.save   v.xunit28-47.vtemp2#branch
.save   v.xunit28-48.vtemp2#branch
.save   v.xunit28-49.vtemp2#branch
.save   v.xunit28-50.vtemp2#branch

.save   v.xunit29-1.vtemp2#branch
.save   v.xunit29-2.vtemp2#branch
.save   v.xunit29-3.vtemp2#branch
.save   v.xunit29-4.vtemp2#branch
.save   v.xunit29-5.vtemp2#branch
.save   v.xunit29-6.vtemp2#branch
.save   v.xunit29-7.vtemp2#branch
.save   v.xunit29-8.vtemp2#branch
.save   v.xunit29-9.vtemp2#branch
.save   v.xunit29-10.vtemp2#branch
.save   v.xunit29-11.vtemp2#branch
.save   v.xunit29-12.vtemp2#branch
.save   v.xunit29-13.vtemp2#branch
.save   v.xunit29-14.vtemp2#branch
.save   v.xunit29-15.vtemp2#branch
.save   v.xunit29-16.vtemp2#branch
.save   v.xunit29-17.vtemp2#branch
.save   v.xunit29-18.vtemp2#branch
.save   v.xunit29-19.vtemp2#branch
.save   v.xunit29-20.vtemp2#branch
.save   v.xunit29-21.vtemp2#branch
.save   v.xunit29-22.vtemp2#branch
.save   v.xunit29-23.vtemp2#branch
.save   v.xunit29-24.vtemp2#branch
.save   v.xunit29-25.vtemp2#branch
.save   v.xunit29-26.vtemp2#branch
.save   v.xunit29-27.vtemp2#branch
.save   v.xunit29-28.vtemp2#branch
.save   v.xunit29-29.vtemp2#branch
.save   v.xunit29-30.vtemp2#branch
.save   v.xunit29-31.vtemp2#branch
.save   v.xunit29-32.vtemp2#branch
.save   v.xunit29-33.vtemp2#branch
.save   v.xunit29-34.vtemp2#branch
.save   v.xunit29-35.vtemp2#branch
.save   v.xunit29-36.vtemp2#branch
.save   v.xunit29-37.vtemp2#branch
.save   v.xunit29-38.vtemp2#branch
.save   v.xunit29-39.vtemp2#branch
.save   v.xunit29-40.vtemp2#branch
.save   v.xunit29-41.vtemp2#branch
.save   v.xunit29-42.vtemp2#branch
.save   v.xunit29-43.vtemp2#branch
.save   v.xunit29-44.vtemp2#branch
.save   v.xunit29-45.vtemp2#branch
.save   v.xunit29-46.vtemp2#branch
.save   v.xunit29-47.vtemp2#branch
.save   v.xunit29-48.vtemp2#branch
.save   v.xunit29-49.vtemp2#branch
.save   v.xunit29-50.vtemp2#branch

.save   v.xunit30-1.vtemp2#branch
.save   v.xunit30-2.vtemp2#branch
.save   v.xunit30-3.vtemp2#branch
.save   v.xunit30-4.vtemp2#branch
.save   v.xunit30-5.vtemp2#branch
.save   v.xunit30-6.vtemp2#branch
.save   v.xunit30-7.vtemp2#branch
.save   v.xunit30-8.vtemp2#branch
.save   v.xunit30-9.vtemp2#branch
.save   v.xunit30-10.vtemp2#branch
.save   v.xunit30-11.vtemp2#branch
.save   v.xunit30-12.vtemp2#branch
.save   v.xunit30-13.vtemp2#branch
.save   v.xunit30-14.vtemp2#branch
.save   v.xunit30-15.vtemp2#branch
.save   v.xunit30-16.vtemp2#branch
.save   v.xunit30-17.vtemp2#branch
.save   v.xunit30-18.vtemp2#branch
.save   v.xunit30-19.vtemp2#branch
.save   v.xunit30-20.vtemp2#branch
.save   v.xunit30-21.vtemp2#branch
.save   v.xunit30-22.vtemp2#branch
.save   v.xunit30-23.vtemp2#branch
.save   v.xunit30-24.vtemp2#branch
.save   v.xunit30-25.vtemp2#branch
.save   v.xunit30-26.vtemp2#branch
.save   v.xunit30-27.vtemp2#branch
.save   v.xunit30-28.vtemp2#branch
.save   v.xunit30-29.vtemp2#branch
.save   v.xunit30-30.vtemp2#branch
.save   v.xunit30-31.vtemp2#branch
.save   v.xunit30-32.vtemp2#branch
.save   v.xunit30-33.vtemp2#branch
.save   v.xunit30-34.vtemp2#branch
.save   v.xunit30-35.vtemp2#branch
.save   v.xunit30-36.vtemp2#branch
.save   v.xunit30-37.vtemp2#branch
.save   v.xunit30-38.vtemp2#branch
.save   v.xunit30-39.vtemp2#branch
.save   v.xunit30-40.vtemp2#branch
.save   v.xunit30-41.vtemp2#branch
.save   v.xunit30-42.vtemp2#branch
.save   v.xunit30-43.vtemp2#branch
.save   v.xunit30-44.vtemp2#branch
.save   v.xunit30-45.vtemp2#branch
.save   v.xunit30-46.vtemp2#branch
.save   v.xunit30-47.vtemp2#branch
.save   v.xunit30-48.vtemp2#branch
.save   v.xunit30-49.vtemp2#branch
.save   v.xunit30-50.vtemp2#branch

.save   v.xunit31-1.vtemp2#branch
.save   v.xunit31-2.vtemp2#branch
.save   v.xunit31-3.vtemp2#branch
.save   v.xunit31-4.vtemp2#branch
.save   v.xunit31-5.vtemp2#branch
.save   v.xunit31-6.vtemp2#branch
.save   v.xunit31-7.vtemp2#branch
.save   v.xunit31-8.vtemp2#branch
.save   v.xunit31-9.vtemp2#branch
.save   v.xunit31-10.vtemp2#branch
.save   v.xunit31-11.vtemp2#branch
.save   v.xunit31-12.vtemp2#branch
.save   v.xunit31-13.vtemp2#branch
.save   v.xunit31-14.vtemp2#branch
.save   v.xunit31-15.vtemp2#branch
.save   v.xunit31-16.vtemp2#branch
.save   v.xunit31-17.vtemp2#branch
.save   v.xunit31-18.vtemp2#branch
.save   v.xunit31-19.vtemp2#branch
.save   v.xunit31-20.vtemp2#branch
.save   v.xunit31-21.vtemp2#branch
.save   v.xunit31-22.vtemp2#branch
.save   v.xunit31-23.vtemp2#branch
.save   v.xunit31-24.vtemp2#branch
.save   v.xunit31-25.vtemp2#branch
.save   v.xunit31-26.vtemp2#branch
.save   v.xunit31-27.vtemp2#branch
.save   v.xunit31-28.vtemp2#branch
.save   v.xunit31-29.vtemp2#branch
.save   v.xunit31-30.vtemp2#branch
.save   v.xunit31-31.vtemp2#branch
.save   v.xunit31-32.vtemp2#branch
.save   v.xunit31-33.vtemp2#branch
.save   v.xunit31-34.vtemp2#branch
.save   v.xunit31-35.vtemp2#branch
.save   v.xunit31-36.vtemp2#branch
.save   v.xunit31-37.vtemp2#branch
.save   v.xunit31-38.vtemp2#branch
.save   v.xunit31-39.vtemp2#branch
.save   v.xunit31-40.vtemp2#branch
.save   v.xunit31-41.vtemp2#branch
.save   v.xunit31-42.vtemp2#branch
.save   v.xunit31-43.vtemp2#branch
.save   v.xunit31-44.vtemp2#branch
.save   v.xunit31-45.vtemp2#branch
.save   v.xunit31-46.vtemp2#branch
.save   v.xunit31-47.vtemp2#branch
.save   v.xunit31-48.vtemp2#branch
.save   v.xunit31-49.vtemp2#branch
.save   v.xunit31-50.vtemp2#branch

.save   v.xunit32-1.vtemp2#branch
.save   v.xunit32-2.vtemp2#branch
.save   v.xunit32-3.vtemp2#branch
.save   v.xunit32-4.vtemp2#branch
.save   v.xunit32-5.vtemp2#branch
.save   v.xunit32-6.vtemp2#branch
.save   v.xunit32-7.vtemp2#branch
.save   v.xunit32-8.vtemp2#branch
.save   v.xunit32-9.vtemp2#branch
.save   v.xunit32-10.vtemp2#branch
.save   v.xunit32-11.vtemp2#branch
.save   v.xunit32-12.vtemp2#branch
.save   v.xunit32-13.vtemp2#branch
.save   v.xunit32-14.vtemp2#branch
.save   v.xunit32-15.vtemp2#branch
.save   v.xunit32-16.vtemp2#branch
.save   v.xunit32-17.vtemp2#branch
.save   v.xunit32-18.vtemp2#branch
.save   v.xunit32-19.vtemp2#branch
.save   v.xunit32-20.vtemp2#branch
.save   v.xunit32-21.vtemp2#branch
.save   v.xunit32-22.vtemp2#branch
.save   v.xunit32-23.vtemp2#branch
.save   v.xunit32-24.vtemp2#branch
.save   v.xunit32-25.vtemp2#branch
.save   v.xunit32-26.vtemp2#branch
.save   v.xunit32-27.vtemp2#branch
.save   v.xunit32-28.vtemp2#branch
.save   v.xunit32-29.vtemp2#branch
.save   v.xunit32-30.vtemp2#branch
.save   v.xunit32-31.vtemp2#branch
.save   v.xunit32-32.vtemp2#branch
.save   v.xunit32-33.vtemp2#branch
.save   v.xunit32-34.vtemp2#branch
.save   v.xunit32-35.vtemp2#branch
.save   v.xunit32-36.vtemp2#branch
.save   v.xunit32-37.vtemp2#branch
.save   v.xunit32-38.vtemp2#branch
.save   v.xunit32-39.vtemp2#branch
.save   v.xunit32-40.vtemp2#branch
.save   v.xunit32-41.vtemp2#branch
.save   v.xunit32-42.vtemp2#branch
.save   v.xunit32-43.vtemp2#branch
.save   v.xunit32-44.vtemp2#branch
.save   v.xunit32-45.vtemp2#branch
.save   v.xunit32-46.vtemp2#branch
.save   v.xunit32-47.vtemp2#branch
.save   v.xunit32-48.vtemp2#branch
.save   v.xunit32-49.vtemp2#branch
.save   v.xunit32-50.vtemp2#branch

.save   v.xunit33-1.vtemp2#branch
.save   v.xunit33-2.vtemp2#branch
.save   v.xunit33-3.vtemp2#branch
.save   v.xunit33-4.vtemp2#branch
.save   v.xunit33-5.vtemp2#branch
.save   v.xunit33-6.vtemp2#branch
.save   v.xunit33-7.vtemp2#branch
.save   v.xunit33-8.vtemp2#branch
.save   v.xunit33-9.vtemp2#branch
.save   v.xunit33-10.vtemp2#branch
.save   v.xunit33-11.vtemp2#branch
.save   v.xunit33-12.vtemp2#branch
.save   v.xunit33-13.vtemp2#branch
.save   v.xunit33-14.vtemp2#branch
.save   v.xunit33-15.vtemp2#branch
.save   v.xunit33-16.vtemp2#branch
.save   v.xunit33-17.vtemp2#branch
.save   v.xunit33-18.vtemp2#branch
.save   v.xunit33-19.vtemp2#branch
.save   v.xunit33-20.vtemp2#branch
.save   v.xunit33-21.vtemp2#branch
.save   v.xunit33-22.vtemp2#branch
.save   v.xunit33-23.vtemp2#branch
.save   v.xunit33-24.vtemp2#branch
.save   v.xunit33-25.vtemp2#branch
.save   v.xunit33-26.vtemp2#branch
.save   v.xunit33-27.vtemp2#branch
.save   v.xunit33-28.vtemp2#branch
.save   v.xunit33-29.vtemp2#branch
.save   v.xunit33-30.vtemp2#branch
.save   v.xunit33-31.vtemp2#branch
.save   v.xunit33-32.vtemp2#branch
.save   v.xunit33-33.vtemp2#branch
.save   v.xunit33-34.vtemp2#branch
.save   v.xunit33-35.vtemp2#branch
.save   v.xunit33-36.vtemp2#branch
.save   v.xunit33-37.vtemp2#branch
.save   v.xunit33-38.vtemp2#branch
.save   v.xunit33-39.vtemp2#branch
.save   v.xunit33-40.vtemp2#branch
.save   v.xunit33-41.vtemp2#branch
.save   v.xunit33-42.vtemp2#branch
.save   v.xunit33-43.vtemp2#branch
.save   v.xunit33-44.vtemp2#branch
.save   v.xunit33-45.vtemp2#branch
.save   v.xunit33-46.vtemp2#branch
.save   v.xunit33-47.vtemp2#branch
.save   v.xunit33-48.vtemp2#branch
.save   v.xunit33-49.vtemp2#branch
.save   v.xunit33-50.vtemp2#branch

.save   v.xunit34-1.vtemp2#branch
.save   v.xunit34-2.vtemp2#branch
.save   v.xunit34-3.vtemp2#branch
.save   v.xunit34-4.vtemp2#branch
.save   v.xunit34-5.vtemp2#branch
.save   v.xunit34-6.vtemp2#branch
.save   v.xunit34-7.vtemp2#branch
.save   v.xunit34-8.vtemp2#branch
.save   v.xunit34-9.vtemp2#branch
.save   v.xunit34-10.vtemp2#branch
.save   v.xunit34-11.vtemp2#branch
.save   v.xunit34-12.vtemp2#branch
.save   v.xunit34-13.vtemp2#branch
.save   v.xunit34-14.vtemp2#branch
.save   v.xunit34-15.vtemp2#branch
.save   v.xunit34-16.vtemp2#branch
.save   v.xunit34-17.vtemp2#branch
.save   v.xunit34-18.vtemp2#branch
.save   v.xunit34-19.vtemp2#branch
.save   v.xunit34-20.vtemp2#branch
.save   v.xunit34-21.vtemp2#branch
.save   v.xunit34-22.vtemp2#branch
.save   v.xunit34-23.vtemp2#branch
.save   v.xunit34-24.vtemp2#branch
.save   v.xunit34-25.vtemp2#branch
.save   v.xunit34-26.vtemp2#branch
.save   v.xunit34-27.vtemp2#branch
.save   v.xunit34-28.vtemp2#branch
.save   v.xunit34-29.vtemp2#branch
.save   v.xunit34-30.vtemp2#branch
.save   v.xunit34-31.vtemp2#branch
.save   v.xunit34-32.vtemp2#branch
.save   v.xunit34-33.vtemp2#branch
.save   v.xunit34-34.vtemp2#branch
.save   v.xunit34-35.vtemp2#branch
.save   v.xunit34-36.vtemp2#branch
.save   v.xunit34-37.vtemp2#branch
.save   v.xunit34-38.vtemp2#branch
.save   v.xunit34-39.vtemp2#branch
.save   v.xunit34-40.vtemp2#branch
.save   v.xunit34-41.vtemp2#branch
.save   v.xunit34-42.vtemp2#branch
.save   v.xunit34-43.vtemp2#branch
.save   v.xunit34-44.vtemp2#branch
.save   v.xunit34-45.vtemp2#branch
.save   v.xunit34-46.vtemp2#branch
.save   v.xunit34-47.vtemp2#branch
.save   v.xunit34-48.vtemp2#branch
.save   v.xunit34-49.vtemp2#branch
.save   v.xunit34-50.vtemp2#branch

.save   v.xunit35-1.vtemp2#branch
.save   v.xunit35-2.vtemp2#branch
.save   v.xunit35-3.vtemp2#branch
.save   v.xunit35-4.vtemp2#branch
.save   v.xunit35-5.vtemp2#branch
.save   v.xunit35-6.vtemp2#branch
.save   v.xunit35-7.vtemp2#branch
.save   v.xunit35-8.vtemp2#branch
.save   v.xunit35-9.vtemp2#branch
.save   v.xunit35-10.vtemp2#branch
.save   v.xunit35-11.vtemp2#branch
.save   v.xunit35-12.vtemp2#branch
.save   v.xunit35-13.vtemp2#branch
.save   v.xunit35-14.vtemp2#branch
.save   v.xunit35-15.vtemp2#branch
.save   v.xunit35-16.vtemp2#branch
.save   v.xunit35-17.vtemp2#branch
.save   v.xunit35-18.vtemp2#branch
.save   v.xunit35-19.vtemp2#branch
.save   v.xunit35-20.vtemp2#branch
.save   v.xunit35-21.vtemp2#branch
.save   v.xunit35-22.vtemp2#branch
.save   v.xunit35-23.vtemp2#branch
.save   v.xunit35-24.vtemp2#branch
.save   v.xunit35-25.vtemp2#branch
.save   v.xunit35-26.vtemp2#branch
.save   v.xunit35-27.vtemp2#branch
.save   v.xunit35-28.vtemp2#branch
.save   v.xunit35-29.vtemp2#branch
.save   v.xunit35-30.vtemp2#branch
.save   v.xunit35-31.vtemp2#branch
.save   v.xunit35-32.vtemp2#branch
.save   v.xunit35-33.vtemp2#branch
.save   v.xunit35-34.vtemp2#branch
.save   v.xunit35-35.vtemp2#branch
.save   v.xunit35-36.vtemp2#branch
.save   v.xunit35-37.vtemp2#branch
.save   v.xunit35-38.vtemp2#branch
.save   v.xunit35-39.vtemp2#branch
.save   v.xunit35-40.vtemp2#branch
.save   v.xunit35-41.vtemp2#branch
.save   v.xunit35-42.vtemp2#branch
.save   v.xunit35-43.vtemp2#branch
.save   v.xunit35-44.vtemp2#branch
.save   v.xunit35-45.vtemp2#branch
.save   v.xunit35-46.vtemp2#branch
.save   v.xunit35-47.vtemp2#branch
.save   v.xunit35-48.vtemp2#branch
.save   v.xunit35-49.vtemp2#branch
.save   v.xunit35-50.vtemp2#branch

.save   v.xunit36-1.vtemp2#branch
.save   v.xunit36-2.vtemp2#branch
.save   v.xunit36-3.vtemp2#branch
.save   v.xunit36-4.vtemp2#branch
.save   v.xunit36-5.vtemp2#branch
.save   v.xunit36-6.vtemp2#branch
.save   v.xunit36-7.vtemp2#branch
.save   v.xunit36-8.vtemp2#branch
.save   v.xunit36-9.vtemp2#branch
.save   v.xunit36-10.vtemp2#branch
.save   v.xunit36-11.vtemp2#branch
.save   v.xunit36-12.vtemp2#branch
.save   v.xunit36-13.vtemp2#branch
.save   v.xunit36-14.vtemp2#branch
.save   v.xunit36-15.vtemp2#branch
.save   v.xunit36-16.vtemp2#branch
.save   v.xunit36-17.vtemp2#branch
.save   v.xunit36-18.vtemp2#branch
.save   v.xunit36-19.vtemp2#branch
.save   v.xunit36-20.vtemp2#branch
.save   v.xunit36-21.vtemp2#branch
.save   v.xunit36-22.vtemp2#branch
.save   v.xunit36-23.vtemp2#branch
.save   v.xunit36-24.vtemp2#branch
.save   v.xunit36-25.vtemp2#branch
.save   v.xunit36-26.vtemp2#branch
.save   v.xunit36-27.vtemp2#branch
.save   v.xunit36-28.vtemp2#branch
.save   v.xunit36-29.vtemp2#branch
.save   v.xunit36-30.vtemp2#branch
.save   v.xunit36-31.vtemp2#branch
.save   v.xunit36-32.vtemp2#branch
.save   v.xunit36-33.vtemp2#branch
.save   v.xunit36-34.vtemp2#branch
.save   v.xunit36-35.vtemp2#branch
.save   v.xunit36-36.vtemp2#branch
.save   v.xunit36-37.vtemp2#branch
.save   v.xunit36-38.vtemp2#branch
.save   v.xunit36-39.vtemp2#branch
.save   v.xunit36-40.vtemp2#branch
.save   v.xunit36-41.vtemp2#branch
.save   v.xunit36-42.vtemp2#branch
.save   v.xunit36-43.vtemp2#branch
.save   v.xunit36-44.vtemp2#branch
.save   v.xunit36-45.vtemp2#branch
.save   v.xunit36-46.vtemp2#branch
.save   v.xunit36-47.vtemp2#branch
.save   v.xunit36-48.vtemp2#branch
.save   v.xunit36-49.vtemp2#branch
.save   v.xunit36-50.vtemp2#branch

.save   v.xunit37-1.vtemp2#branch
.save   v.xunit37-2.vtemp2#branch
.save   v.xunit37-3.vtemp2#branch
.save   v.xunit37-4.vtemp2#branch
.save   v.xunit37-5.vtemp2#branch
.save   v.xunit37-6.vtemp2#branch
.save   v.xunit37-7.vtemp2#branch
.save   v.xunit37-8.vtemp2#branch
.save   v.xunit37-9.vtemp2#branch
.save   v.xunit37-10.vtemp2#branch
.save   v.xunit37-11.vtemp2#branch
.save   v.xunit37-12.vtemp2#branch
.save   v.xunit37-13.vtemp2#branch
.save   v.xunit37-14.vtemp2#branch
.save   v.xunit37-15.vtemp2#branch
.save   v.xunit37-16.vtemp2#branch
.save   v.xunit37-17.vtemp2#branch
.save   v.xunit37-18.vtemp2#branch
.save   v.xunit37-19.vtemp2#branch
.save   v.xunit37-20.vtemp2#branch
.save   v.xunit37-21.vtemp2#branch
.save   v.xunit37-22.vtemp2#branch
.save   v.xunit37-23.vtemp2#branch
.save   v.xunit37-24.vtemp2#branch
.save   v.xunit37-25.vtemp2#branch
.save   v.xunit37-26.vtemp2#branch
.save   v.xunit37-27.vtemp2#branch
.save   v.xunit37-28.vtemp2#branch
.save   v.xunit37-29.vtemp2#branch
.save   v.xunit37-30.vtemp2#branch
.save   v.xunit37-31.vtemp2#branch
.save   v.xunit37-32.vtemp2#branch
.save   v.xunit37-33.vtemp2#branch
.save   v.xunit37-34.vtemp2#branch
.save   v.xunit37-35.vtemp2#branch
.save   v.xunit37-36.vtemp2#branch
.save   v.xunit37-37.vtemp2#branch
.save   v.xunit37-38.vtemp2#branch
.save   v.xunit37-39.vtemp2#branch
.save   v.xunit37-40.vtemp2#branch
.save   v.xunit37-41.vtemp2#branch
.save   v.xunit37-42.vtemp2#branch
.save   v.xunit37-43.vtemp2#branch
.save   v.xunit37-44.vtemp2#branch
.save   v.xunit37-45.vtemp2#branch
.save   v.xunit37-46.vtemp2#branch
.save   v.xunit37-47.vtemp2#branch
.save   v.xunit37-48.vtemp2#branch
.save   v.xunit37-49.vtemp2#branch
.save   v.xunit37-50.vtemp2#branch

.save   v.xunit38-1.vtemp2#branch
.save   v.xunit38-2.vtemp2#branch
.save   v.xunit38-3.vtemp2#branch
.save   v.xunit38-4.vtemp2#branch
.save   v.xunit38-5.vtemp2#branch
.save   v.xunit38-6.vtemp2#branch
.save   v.xunit38-7.vtemp2#branch
.save   v.xunit38-8.vtemp2#branch
.save   v.xunit38-9.vtemp2#branch
.save   v.xunit38-10.vtemp2#branch
.save   v.xunit38-11.vtemp2#branch
.save   v.xunit38-12.vtemp2#branch
.save   v.xunit38-13.vtemp2#branch
.save   v.xunit38-14.vtemp2#branch
.save   v.xunit38-15.vtemp2#branch
.save   v.xunit38-16.vtemp2#branch
.save   v.xunit38-17.vtemp2#branch
.save   v.xunit38-18.vtemp2#branch
.save   v.xunit38-19.vtemp2#branch
.save   v.xunit38-20.vtemp2#branch
.save   v.xunit38-21.vtemp2#branch
.save   v.xunit38-22.vtemp2#branch
.save   v.xunit38-23.vtemp2#branch
.save   v.xunit38-24.vtemp2#branch
.save   v.xunit38-25.vtemp2#branch
.save   v.xunit38-26.vtemp2#branch
.save   v.xunit38-27.vtemp2#branch
.save   v.xunit38-28.vtemp2#branch
.save   v.xunit38-29.vtemp2#branch
.save   v.xunit38-30.vtemp2#branch
.save   v.xunit38-31.vtemp2#branch
.save   v.xunit38-32.vtemp2#branch
.save   v.xunit38-33.vtemp2#branch
.save   v.xunit38-34.vtemp2#branch
.save   v.xunit38-35.vtemp2#branch
.save   v.xunit38-36.vtemp2#branch
.save   v.xunit38-37.vtemp2#branch
.save   v.xunit38-38.vtemp2#branch
.save   v.xunit38-39.vtemp2#branch
.save   v.xunit38-40.vtemp2#branch
.save   v.xunit38-41.vtemp2#branch
.save   v.xunit38-42.vtemp2#branch
.save   v.xunit38-43.vtemp2#branch
.save   v.xunit38-44.vtemp2#branch
.save   v.xunit38-45.vtemp2#branch
.save   v.xunit38-46.vtemp2#branch
.save   v.xunit38-47.vtemp2#branch
.save   v.xunit38-48.vtemp2#branch
.save   v.xunit38-49.vtemp2#branch
.save   v.xunit38-50.vtemp2#branch

.save   v.xunit39-1.vtemp2#branch
.save   v.xunit39-2.vtemp2#branch
.save   v.xunit39-3.vtemp2#branch
.save   v.xunit39-4.vtemp2#branch
.save   v.xunit39-5.vtemp2#branch
.save   v.xunit39-6.vtemp2#branch
.save   v.xunit39-7.vtemp2#branch
.save   v.xunit39-8.vtemp2#branch
.save   v.xunit39-9.vtemp2#branch
.save   v.xunit39-10.vtemp2#branch
.save   v.xunit39-11.vtemp2#branch
.save   v.xunit39-12.vtemp2#branch
.save   v.xunit39-13.vtemp2#branch
.save   v.xunit39-14.vtemp2#branch
.save   v.xunit39-15.vtemp2#branch
.save   v.xunit39-16.vtemp2#branch
.save   v.xunit39-17.vtemp2#branch
.save   v.xunit39-18.vtemp2#branch
.save   v.xunit39-19.vtemp2#branch
.save   v.xunit39-20.vtemp2#branch
.save   v.xunit39-21.vtemp2#branch
.save   v.xunit39-22.vtemp2#branch
.save   v.xunit39-23.vtemp2#branch
.save   v.xunit39-24.vtemp2#branch
.save   v.xunit39-25.vtemp2#branch
.save   v.xunit39-26.vtemp2#branch
.save   v.xunit39-27.vtemp2#branch
.save   v.xunit39-28.vtemp2#branch
.save   v.xunit39-29.vtemp2#branch
.save   v.xunit39-30.vtemp2#branch
.save   v.xunit39-31.vtemp2#branch
.save   v.xunit39-32.vtemp2#branch
.save   v.xunit39-33.vtemp2#branch
.save   v.xunit39-34.vtemp2#branch
.save   v.xunit39-35.vtemp2#branch
.save   v.xunit39-36.vtemp2#branch
.save   v.xunit39-37.vtemp2#branch
.save   v.xunit39-38.vtemp2#branch
.save   v.xunit39-39.vtemp2#branch
.save   v.xunit39-40.vtemp2#branch
.save   v.xunit39-41.vtemp2#branch
.save   v.xunit39-42.vtemp2#branch
.save   v.xunit39-43.vtemp2#branch
.save   v.xunit39-44.vtemp2#branch
.save   v.xunit39-45.vtemp2#branch
.save   v.xunit39-46.vtemp2#branch
.save   v.xunit39-47.vtemp2#branch
.save   v.xunit39-48.vtemp2#branch
.save   v.xunit39-49.vtemp2#branch
.save   v.xunit39-50.vtemp2#branch

.save   v.xunit40-1.vtemp2#branch
.save   v.xunit40-2.vtemp2#branch
.save   v.xunit40-3.vtemp2#branch
.save   v.xunit40-4.vtemp2#branch
.save   v.xunit40-5.vtemp2#branch
.save   v.xunit40-6.vtemp2#branch
.save   v.xunit40-7.vtemp2#branch
.save   v.xunit40-8.vtemp2#branch
.save   v.xunit40-9.vtemp2#branch
.save   v.xunit40-10.vtemp2#branch
.save   v.xunit40-11.vtemp2#branch
.save   v.xunit40-12.vtemp2#branch
.save   v.xunit40-13.vtemp2#branch
.save   v.xunit40-14.vtemp2#branch
.save   v.xunit40-15.vtemp2#branch
.save   v.xunit40-16.vtemp2#branch
.save   v.xunit40-17.vtemp2#branch
.save   v.xunit40-18.vtemp2#branch
.save   v.xunit40-19.vtemp2#branch
.save   v.xunit40-20.vtemp2#branch
.save   v.xunit40-21.vtemp2#branch
.save   v.xunit40-22.vtemp2#branch
.save   v.xunit40-23.vtemp2#branch
.save   v.xunit40-24.vtemp2#branch
.save   v.xunit40-25.vtemp2#branch
.save   v.xunit40-26.vtemp2#branch
.save   v.xunit40-27.vtemp2#branch
.save   v.xunit40-28.vtemp2#branch
.save   v.xunit40-29.vtemp2#branch
.save   v.xunit40-30.vtemp2#branch
.save   v.xunit40-31.vtemp2#branch
.save   v.xunit40-32.vtemp2#branch
.save   v.xunit40-33.vtemp2#branch
.save   v.xunit40-34.vtemp2#branch
.save   v.xunit40-35.vtemp2#branch
.save   v.xunit40-36.vtemp2#branch
.save   v.xunit40-37.vtemp2#branch
.save   v.xunit40-38.vtemp2#branch
.save   v.xunit40-39.vtemp2#branch
.save   v.xunit40-40.vtemp2#branch
.save   v.xunit40-41.vtemp2#branch
.save   v.xunit40-42.vtemp2#branch
.save   v.xunit40-43.vtemp2#branch
.save   v.xunit40-44.vtemp2#branch
.save   v.xunit40-45.vtemp2#branch
.save   v.xunit40-46.vtemp2#branch
.save   v.xunit40-47.vtemp2#branch
.save   v.xunit40-48.vtemp2#branch
.save   v.xunit40-49.vtemp2#branch
.save   v.xunit40-50.vtemp2#branch

.save   v.xunit41-1.vtemp2#branch
.save   v.xunit41-2.vtemp2#branch
.save   v.xunit41-3.vtemp2#branch
.save   v.xunit41-4.vtemp2#branch
.save   v.xunit41-5.vtemp2#branch
.save   v.xunit41-6.vtemp2#branch
.save   v.xunit41-7.vtemp2#branch
.save   v.xunit41-8.vtemp2#branch
.save   v.xunit41-9.vtemp2#branch
.save   v.xunit41-10.vtemp2#branch
.save   v.xunit41-11.vtemp2#branch
.save   v.xunit41-12.vtemp2#branch
.save   v.xunit41-13.vtemp2#branch
.save   v.xunit41-14.vtemp2#branch
.save   v.xunit41-15.vtemp2#branch
.save   v.xunit41-16.vtemp2#branch
.save   v.xunit41-17.vtemp2#branch
.save   v.xunit41-18.vtemp2#branch
.save   v.xunit41-19.vtemp2#branch
.save   v.xunit41-20.vtemp2#branch
.save   v.xunit41-21.vtemp2#branch
.save   v.xunit41-22.vtemp2#branch
.save   v.xunit41-23.vtemp2#branch
.save   v.xunit41-24.vtemp2#branch
.save   v.xunit41-25.vtemp2#branch
.save   v.xunit41-26.vtemp2#branch
.save   v.xunit41-27.vtemp2#branch
.save   v.xunit41-28.vtemp2#branch
.save   v.xunit41-29.vtemp2#branch
.save   v.xunit41-30.vtemp2#branch
.save   v.xunit41-31.vtemp2#branch
.save   v.xunit41-32.vtemp2#branch
.save   v.xunit41-33.vtemp2#branch
.save   v.xunit41-34.vtemp2#branch
.save   v.xunit41-35.vtemp2#branch
.save   v.xunit41-36.vtemp2#branch
.save   v.xunit41-37.vtemp2#branch
.save   v.xunit41-38.vtemp2#branch
.save   v.xunit41-39.vtemp2#branch
.save   v.xunit41-40.vtemp2#branch
.save   v.xunit41-41.vtemp2#branch
.save   v.xunit41-42.vtemp2#branch
.save   v.xunit41-43.vtemp2#branch
.save   v.xunit41-44.vtemp2#branch
.save   v.xunit41-45.vtemp2#branch
.save   v.xunit41-46.vtemp2#branch
.save   v.xunit41-47.vtemp2#branch
.save   v.xunit41-48.vtemp2#branch
.save   v.xunit41-49.vtemp2#branch
.save   v.xunit41-50.vtemp2#branch

.save   v.xunit42-1.vtemp2#branch
.save   v.xunit42-2.vtemp2#branch
.save   v.xunit42-3.vtemp2#branch
.save   v.xunit42-4.vtemp2#branch
.save   v.xunit42-5.vtemp2#branch
.save   v.xunit42-6.vtemp2#branch
.save   v.xunit42-7.vtemp2#branch
.save   v.xunit42-8.vtemp2#branch
.save   v.xunit42-9.vtemp2#branch
.save   v.xunit42-10.vtemp2#branch
.save   v.xunit42-11.vtemp2#branch
.save   v.xunit42-12.vtemp2#branch
.save   v.xunit42-13.vtemp2#branch
.save   v.xunit42-14.vtemp2#branch
.save   v.xunit42-15.vtemp2#branch
.save   v.xunit42-16.vtemp2#branch
.save   v.xunit42-17.vtemp2#branch
.save   v.xunit42-18.vtemp2#branch
.save   v.xunit42-19.vtemp2#branch
.save   v.xunit42-20.vtemp2#branch
.save   v.xunit42-21.vtemp2#branch
.save   v.xunit42-22.vtemp2#branch
.save   v.xunit42-23.vtemp2#branch
.save   v.xunit42-24.vtemp2#branch
.save   v.xunit42-25.vtemp2#branch
.save   v.xunit42-26.vtemp2#branch
.save   v.xunit42-27.vtemp2#branch
.save   v.xunit42-28.vtemp2#branch
.save   v.xunit42-29.vtemp2#branch
.save   v.xunit42-30.vtemp2#branch
.save   v.xunit42-31.vtemp2#branch
.save   v.xunit42-32.vtemp2#branch
.save   v.xunit42-33.vtemp2#branch
.save   v.xunit42-34.vtemp2#branch
.save   v.xunit42-35.vtemp2#branch
.save   v.xunit42-36.vtemp2#branch
.save   v.xunit42-37.vtemp2#branch
.save   v.xunit42-38.vtemp2#branch
.save   v.xunit42-39.vtemp2#branch
.save   v.xunit42-40.vtemp2#branch
.save   v.xunit42-41.vtemp2#branch
.save   v.xunit42-42.vtemp2#branch
.save   v.xunit42-43.vtemp2#branch
.save   v.xunit42-44.vtemp2#branch
.save   v.xunit42-45.vtemp2#branch
.save   v.xunit42-46.vtemp2#branch
.save   v.xunit42-47.vtemp2#branch
.save   v.xunit42-48.vtemp2#branch
.save   v.xunit42-49.vtemp2#branch
.save   v.xunit42-50.vtemp2#branch

.save   v.xunit43-1.vtemp2#branch
.save   v.xunit43-2.vtemp2#branch
.save   v.xunit43-3.vtemp2#branch
.save   v.xunit43-4.vtemp2#branch
.save   v.xunit43-5.vtemp2#branch
.save   v.xunit43-6.vtemp2#branch
.save   v.xunit43-7.vtemp2#branch
.save   v.xunit43-8.vtemp2#branch
.save   v.xunit43-9.vtemp2#branch
.save   v.xunit43-10.vtemp2#branch
.save   v.xunit43-11.vtemp2#branch
.save   v.xunit43-12.vtemp2#branch
.save   v.xunit43-13.vtemp2#branch
.save   v.xunit43-14.vtemp2#branch
.save   v.xunit43-15.vtemp2#branch
.save   v.xunit43-16.vtemp2#branch
.save   v.xunit43-17.vtemp2#branch
.save   v.xunit43-18.vtemp2#branch
.save   v.xunit43-19.vtemp2#branch
.save   v.xunit43-20.vtemp2#branch
.save   v.xunit43-21.vtemp2#branch
.save   v.xunit43-22.vtemp2#branch
.save   v.xunit43-23.vtemp2#branch
.save   v.xunit43-24.vtemp2#branch
.save   v.xunit43-25.vtemp2#branch
.save   v.xunit43-26.vtemp2#branch
.save   v.xunit43-27.vtemp2#branch
.save   v.xunit43-28.vtemp2#branch
.save   v.xunit43-29.vtemp2#branch
.save   v.xunit43-30.vtemp2#branch
.save   v.xunit43-31.vtemp2#branch
.save   v.xunit43-32.vtemp2#branch
.save   v.xunit43-33.vtemp2#branch
.save   v.xunit43-34.vtemp2#branch
.save   v.xunit43-35.vtemp2#branch
.save   v.xunit43-36.vtemp2#branch
.save   v.xunit43-37.vtemp2#branch
.save   v.xunit43-38.vtemp2#branch
.save   v.xunit43-39.vtemp2#branch
.save   v.xunit43-40.vtemp2#branch
.save   v.xunit43-41.vtemp2#branch
.save   v.xunit43-42.vtemp2#branch
.save   v.xunit43-43.vtemp2#branch
.save   v.xunit43-44.vtemp2#branch
.save   v.xunit43-45.vtemp2#branch
.save   v.xunit43-46.vtemp2#branch
.save   v.xunit43-47.vtemp2#branch
.save   v.xunit43-48.vtemp2#branch
.save   v.xunit43-49.vtemp2#branch
.save   v.xunit43-50.vtemp2#branch

.save   v.xunit44-1.vtemp2#branch
.save   v.xunit44-2.vtemp2#branch
.save   v.xunit44-3.vtemp2#branch
.save   v.xunit44-4.vtemp2#branch
.save   v.xunit44-5.vtemp2#branch
.save   v.xunit44-6.vtemp2#branch
.save   v.xunit44-7.vtemp2#branch
.save   v.xunit44-8.vtemp2#branch
.save   v.xunit44-9.vtemp2#branch
.save   v.xunit44-10.vtemp2#branch
.save   v.xunit44-11.vtemp2#branch
.save   v.xunit44-12.vtemp2#branch
.save   v.xunit44-13.vtemp2#branch
.save   v.xunit44-14.vtemp2#branch
.save   v.xunit44-15.vtemp2#branch
.save   v.xunit44-16.vtemp2#branch
.save   v.xunit44-17.vtemp2#branch
.save   v.xunit44-18.vtemp2#branch
.save   v.xunit44-19.vtemp2#branch
.save   v.xunit44-20.vtemp2#branch
.save   v.xunit44-21.vtemp2#branch
.save   v.xunit44-22.vtemp2#branch
.save   v.xunit44-23.vtemp2#branch
.save   v.xunit44-24.vtemp2#branch
.save   v.xunit44-25.vtemp2#branch
.save   v.xunit44-26.vtemp2#branch
.save   v.xunit44-27.vtemp2#branch
.save   v.xunit44-28.vtemp2#branch
.save   v.xunit44-29.vtemp2#branch
.save   v.xunit44-30.vtemp2#branch
.save   v.xunit44-31.vtemp2#branch
.save   v.xunit44-32.vtemp2#branch
.save   v.xunit44-33.vtemp2#branch
.save   v.xunit44-34.vtemp2#branch
.save   v.xunit44-35.vtemp2#branch
.save   v.xunit44-36.vtemp2#branch
.save   v.xunit44-37.vtemp2#branch
.save   v.xunit44-38.vtemp2#branch
.save   v.xunit44-39.vtemp2#branch
.save   v.xunit44-40.vtemp2#branch
.save   v.xunit44-41.vtemp2#branch
.save   v.xunit44-42.vtemp2#branch
.save   v.xunit44-43.vtemp2#branch
.save   v.xunit44-44.vtemp2#branch
.save   v.xunit44-45.vtemp2#branch
.save   v.xunit44-46.vtemp2#branch
.save   v.xunit44-47.vtemp2#branch
.save   v.xunit44-48.vtemp2#branch
.save   v.xunit44-49.vtemp2#branch
.save   v.xunit44-50.vtemp2#branch

.save   v.xunit45-1.vtemp2#branch
.save   v.xunit45-2.vtemp2#branch
.save   v.xunit45-3.vtemp2#branch
.save   v.xunit45-4.vtemp2#branch
.save   v.xunit45-5.vtemp2#branch
.save   v.xunit45-6.vtemp2#branch
.save   v.xunit45-7.vtemp2#branch
.save   v.xunit45-8.vtemp2#branch
.save   v.xunit45-9.vtemp2#branch
.save   v.xunit45-10.vtemp2#branch
.save   v.xunit45-11.vtemp2#branch
.save   v.xunit45-12.vtemp2#branch
.save   v.xunit45-13.vtemp2#branch
.save   v.xunit45-14.vtemp2#branch
.save   v.xunit45-15.vtemp2#branch
.save   v.xunit45-16.vtemp2#branch
.save   v.xunit45-17.vtemp2#branch
.save   v.xunit45-18.vtemp2#branch
.save   v.xunit45-19.vtemp2#branch
.save   v.xunit45-20.vtemp2#branch
.save   v.xunit45-21.vtemp2#branch
.save   v.xunit45-22.vtemp2#branch
.save   v.xunit45-23.vtemp2#branch
.save   v.xunit45-24.vtemp2#branch
.save   v.xunit45-25.vtemp2#branch
.save   v.xunit45-26.vtemp2#branch
.save   v.xunit45-27.vtemp2#branch
.save   v.xunit45-28.vtemp2#branch
.save   v.xunit45-29.vtemp2#branch
.save   v.xunit45-30.vtemp2#branch
.save   v.xunit45-31.vtemp2#branch
.save   v.xunit45-32.vtemp2#branch
.save   v.xunit45-33.vtemp2#branch
.save   v.xunit45-34.vtemp2#branch
.save   v.xunit45-35.vtemp2#branch
.save   v.xunit45-36.vtemp2#branch
.save   v.xunit45-37.vtemp2#branch
.save   v.xunit45-38.vtemp2#branch
.save   v.xunit45-39.vtemp2#branch
.save   v.xunit45-40.vtemp2#branch
.save   v.xunit45-41.vtemp2#branch
.save   v.xunit45-42.vtemp2#branch
.save   v.xunit45-43.vtemp2#branch
.save   v.xunit45-44.vtemp2#branch
.save   v.xunit45-45.vtemp2#branch
.save   v.xunit45-46.vtemp2#branch
.save   v.xunit45-47.vtemp2#branch
.save   v.xunit45-48.vtemp2#branch
.save   v.xunit45-49.vtemp2#branch
.save   v.xunit45-50.vtemp2#branch

.save   v.xunit46-1.vtemp2#branch
.save   v.xunit46-2.vtemp2#branch
.save   v.xunit46-3.vtemp2#branch
.save   v.xunit46-4.vtemp2#branch
.save   v.xunit46-5.vtemp2#branch
.save   v.xunit46-6.vtemp2#branch
.save   v.xunit46-7.vtemp2#branch
.save   v.xunit46-8.vtemp2#branch
.save   v.xunit46-9.vtemp2#branch
.save   v.xunit46-10.vtemp2#branch
.save   v.xunit46-11.vtemp2#branch
.save   v.xunit46-12.vtemp2#branch
.save   v.xunit46-13.vtemp2#branch
.save   v.xunit46-14.vtemp2#branch
.save   v.xunit46-15.vtemp2#branch
.save   v.xunit46-16.vtemp2#branch
.save   v.xunit46-17.vtemp2#branch
.save   v.xunit46-18.vtemp2#branch
.save   v.xunit46-19.vtemp2#branch
.save   v.xunit46-20.vtemp2#branch
.save   v.xunit46-21.vtemp2#branch
.save   v.xunit46-22.vtemp2#branch
.save   v.xunit46-23.vtemp2#branch
.save   v.xunit46-24.vtemp2#branch
.save   v.xunit46-25.vtemp2#branch
.save   v.xunit46-26.vtemp2#branch
.save   v.xunit46-27.vtemp2#branch
.save   v.xunit46-28.vtemp2#branch
.save   v.xunit46-29.vtemp2#branch
.save   v.xunit46-30.vtemp2#branch
.save   v.xunit46-31.vtemp2#branch
.save   v.xunit46-32.vtemp2#branch
.save   v.xunit46-33.vtemp2#branch
.save   v.xunit46-34.vtemp2#branch
.save   v.xunit46-35.vtemp2#branch
.save   v.xunit46-36.vtemp2#branch
.save   v.xunit46-37.vtemp2#branch
.save   v.xunit46-38.vtemp2#branch
.save   v.xunit46-39.vtemp2#branch
.save   v.xunit46-40.vtemp2#branch
.save   v.xunit46-41.vtemp2#branch
.save   v.xunit46-42.vtemp2#branch
.save   v.xunit46-43.vtemp2#branch
.save   v.xunit46-44.vtemp2#branch
.save   v.xunit46-45.vtemp2#branch
.save   v.xunit46-46.vtemp2#branch
.save   v.xunit46-47.vtemp2#branch
.save   v.xunit46-48.vtemp2#branch
.save   v.xunit46-49.vtemp2#branch
.save   v.xunit46-50.vtemp2#branch

.save   v.xunit47-1.vtemp2#branch
.save   v.xunit47-2.vtemp2#branch
.save   v.xunit47-3.vtemp2#branch
.save   v.xunit47-4.vtemp2#branch
.save   v.xunit47-5.vtemp2#branch
.save   v.xunit47-6.vtemp2#branch
.save   v.xunit47-7.vtemp2#branch
.save   v.xunit47-8.vtemp2#branch
.save   v.xunit47-9.vtemp2#branch
.save   v.xunit47-10.vtemp2#branch
.save   v.xunit47-11.vtemp2#branch
.save   v.xunit47-12.vtemp2#branch
.save   v.xunit47-13.vtemp2#branch
.save   v.xunit47-14.vtemp2#branch
.save   v.xunit47-15.vtemp2#branch
.save   v.xunit47-16.vtemp2#branch
.save   v.xunit47-17.vtemp2#branch
.save   v.xunit47-18.vtemp2#branch
.save   v.xunit47-19.vtemp2#branch
.save   v.xunit47-20.vtemp2#branch
.save   v.xunit47-21.vtemp2#branch
.save   v.xunit47-22.vtemp2#branch
.save   v.xunit47-23.vtemp2#branch
.save   v.xunit47-24.vtemp2#branch
.save   v.xunit47-25.vtemp2#branch
.save   v.xunit47-26.vtemp2#branch
.save   v.xunit47-27.vtemp2#branch
.save   v.xunit47-28.vtemp2#branch
.save   v.xunit47-29.vtemp2#branch
.save   v.xunit47-30.vtemp2#branch
.save   v.xunit47-31.vtemp2#branch
.save   v.xunit47-32.vtemp2#branch
.save   v.xunit47-33.vtemp2#branch
.save   v.xunit47-34.vtemp2#branch
.save   v.xunit47-35.vtemp2#branch
.save   v.xunit47-36.vtemp2#branch
.save   v.xunit47-37.vtemp2#branch
.save   v.xunit47-38.vtemp2#branch
.save   v.xunit47-39.vtemp2#branch
.save   v.xunit47-40.vtemp2#branch
.save   v.xunit47-41.vtemp2#branch
.save   v.xunit47-42.vtemp2#branch
.save   v.xunit47-43.vtemp2#branch
.save   v.xunit47-44.vtemp2#branch
.save   v.xunit47-45.vtemp2#branch
.save   v.xunit47-46.vtemp2#branch
.save   v.xunit47-47.vtemp2#branch
.save   v.xunit47-48.vtemp2#branch
.save   v.xunit47-49.vtemp2#branch
.save   v.xunit47-50.vtemp2#branch

.save   v.xunit48-1.vtemp2#branch
.save   v.xunit48-2.vtemp2#branch
.save   v.xunit48-3.vtemp2#branch
.save   v.xunit48-4.vtemp2#branch
.save   v.xunit48-5.vtemp2#branch
.save   v.xunit48-6.vtemp2#branch
.save   v.xunit48-7.vtemp2#branch
.save   v.xunit48-8.vtemp2#branch
.save   v.xunit48-9.vtemp2#branch
.save   v.xunit48-10.vtemp2#branch
.save   v.xunit48-11.vtemp2#branch
.save   v.xunit48-12.vtemp2#branch
.save   v.xunit48-13.vtemp2#branch
.save   v.xunit48-14.vtemp2#branch
.save   v.xunit48-15.vtemp2#branch
.save   v.xunit48-16.vtemp2#branch
.save   v.xunit48-17.vtemp2#branch
.save   v.xunit48-18.vtemp2#branch
.save   v.xunit48-19.vtemp2#branch
.save   v.xunit48-20.vtemp2#branch
.save   v.xunit48-21.vtemp2#branch
.save   v.xunit48-22.vtemp2#branch
.save   v.xunit48-23.vtemp2#branch
.save   v.xunit48-24.vtemp2#branch
.save   v.xunit48-25.vtemp2#branch
.save   v.xunit48-26.vtemp2#branch
.save   v.xunit48-27.vtemp2#branch
.save   v.xunit48-28.vtemp2#branch
.save   v.xunit48-29.vtemp2#branch
.save   v.xunit48-30.vtemp2#branch
.save   v.xunit48-31.vtemp2#branch
.save   v.xunit48-32.vtemp2#branch
.save   v.xunit48-33.vtemp2#branch
.save   v.xunit48-34.vtemp2#branch
.save   v.xunit48-35.vtemp2#branch
.save   v.xunit48-36.vtemp2#branch
.save   v.xunit48-37.vtemp2#branch
.save   v.xunit48-38.vtemp2#branch
.save   v.xunit48-39.vtemp2#branch
.save   v.xunit48-40.vtemp2#branch
.save   v.xunit48-41.vtemp2#branch
.save   v.xunit48-42.vtemp2#branch
.save   v.xunit48-43.vtemp2#branch
.save   v.xunit48-44.vtemp2#branch
.save   v.xunit48-45.vtemp2#branch
.save   v.xunit48-46.vtemp2#branch
.save   v.xunit48-47.vtemp2#branch
.save   v.xunit48-48.vtemp2#branch
.save   v.xunit48-49.vtemp2#branch
.save   v.xunit48-50.vtemp2#branch

.save   v.xunit49-1.vtemp2#branch
.save   v.xunit49-2.vtemp2#branch
.save   v.xunit49-3.vtemp2#branch
.save   v.xunit49-4.vtemp2#branch
.save   v.xunit49-5.vtemp2#branch
.save   v.xunit49-6.vtemp2#branch
.save   v.xunit49-7.vtemp2#branch
.save   v.xunit49-8.vtemp2#branch
.save   v.xunit49-9.vtemp2#branch
.save   v.xunit49-10.vtemp2#branch
.save   v.xunit49-11.vtemp2#branch
.save   v.xunit49-12.vtemp2#branch
.save   v.xunit49-13.vtemp2#branch
.save   v.xunit49-14.vtemp2#branch
.save   v.xunit49-15.vtemp2#branch
.save   v.xunit49-16.vtemp2#branch
.save   v.xunit49-17.vtemp2#branch
.save   v.xunit49-18.vtemp2#branch
.save   v.xunit49-19.vtemp2#branch
.save   v.xunit49-20.vtemp2#branch
.save   v.xunit49-21.vtemp2#branch
.save   v.xunit49-22.vtemp2#branch
.save   v.xunit49-23.vtemp2#branch
.save   v.xunit49-24.vtemp2#branch
.save   v.xunit49-25.vtemp2#branch
.save   v.xunit49-26.vtemp2#branch
.save   v.xunit49-27.vtemp2#branch
.save   v.xunit49-28.vtemp2#branch
.save   v.xunit49-29.vtemp2#branch
.save   v.xunit49-30.vtemp2#branch
.save   v.xunit49-31.vtemp2#branch
.save   v.xunit49-32.vtemp2#branch
.save   v.xunit49-33.vtemp2#branch
.save   v.xunit49-34.vtemp2#branch
.save   v.xunit49-35.vtemp2#branch
.save   v.xunit49-36.vtemp2#branch
.save   v.xunit49-37.vtemp2#branch
.save   v.xunit49-38.vtemp2#branch
.save   v.xunit49-39.vtemp2#branch
.save   v.xunit49-40.vtemp2#branch
.save   v.xunit49-41.vtemp2#branch
.save   v.xunit49-42.vtemp2#branch
.save   v.xunit49-43.vtemp2#branch
.save   v.xunit49-44.vtemp2#branch
.save   v.xunit49-45.vtemp2#branch
.save   v.xunit49-46.vtemp2#branch
.save   v.xunit49-47.vtemp2#branch
.save   v.xunit49-48.vtemp2#branch
.save   v.xunit49-49.vtemp2#branch
.save   v.xunit49-50.vtemp2#branch

.save   v.xunit50-1.vtemp2#branch
.save   v.xunit50-2.vtemp2#branch
.save   v.xunit50-3.vtemp2#branch
.save   v.xunit50-4.vtemp2#branch
.save   v.xunit50-5.vtemp2#branch
.save   v.xunit50-6.vtemp2#branch
.save   v.xunit50-7.vtemp2#branch
.save   v.xunit50-8.vtemp2#branch
.save   v.xunit50-9.vtemp2#branch
.save   v.xunit50-10.vtemp2#branch
.save   v.xunit50-11.vtemp2#branch
.save   v.xunit50-12.vtemp2#branch
.save   v.xunit50-13.vtemp2#branch
.save   v.xunit50-14.vtemp2#branch
.save   v.xunit50-15.vtemp2#branch
.save   v.xunit50-16.vtemp2#branch
.save   v.xunit50-17.vtemp2#branch
.save   v.xunit50-18.vtemp2#branch
.save   v.xunit50-19.vtemp2#branch
.save   v.xunit50-20.vtemp2#branch
.save   v.xunit50-21.vtemp2#branch
.save   v.xunit50-22.vtemp2#branch
.save   v.xunit50-23.vtemp2#branch
.save   v.xunit50-24.vtemp2#branch
.save   v.xunit50-25.vtemp2#branch
.save   v.xunit50-26.vtemp2#branch
.save   v.xunit50-27.vtemp2#branch
.save   v.xunit50-28.vtemp2#branch
.save   v.xunit50-29.vtemp2#branch
.save   v.xunit50-30.vtemp2#branch
.save   v.xunit50-31.vtemp2#branch
.save   v.xunit50-32.vtemp2#branch
.save   v.xunit50-33.vtemp2#branch
.save   v.xunit50-34.vtemp2#branch
.save   v.xunit50-35.vtemp2#branch
.save   v.xunit50-36.vtemp2#branch
.save   v.xunit50-37.vtemp2#branch
.save   v.xunit50-38.vtemp2#branch
.save   v.xunit50-39.vtemp2#branch
.save   v.xunit50-40.vtemp2#branch
.save   v.xunit50-41.vtemp2#branch
.save   v.xunit50-42.vtemp2#branch
.save   v.xunit50-43.vtemp2#branch
.save   v.xunit50-44.vtemp2#branch
.save   v.xunit50-45.vtemp2#branch
.save   v.xunit50-46.vtemp2#branch
.save   v.xunit50-47.vtemp2#branch
.save   v.xunit50-48.vtemp2#branch
.save   v.xunit50-49.vtemp2#branch
.save   v.xunit50-50.vtemp2#branch


.save v(vt1)

.control
set xtrtol=1
let deltime = stime/899
tran $&deltime $&stime uic
linearize
run
write rawfile.raw
set color0=white
set color1=black
set xbrushwidth=2
.endc